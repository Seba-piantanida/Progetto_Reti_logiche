
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 34968; -- 5 + 3 + 20 + 7   (RST) + (CH2-MEM[1]) + 20 CYCLES + (CH1-MEM[6])
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & 
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" ;

    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & 
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" ;

    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & 
		"011010010001101111" &
		"00000000000000000000" &
		"101011000110111000" &
		"00000000000000000000" &
		"0010111110001111" &
		"00000000000000000000" &
		"111101110001111101" &
		"00000000000000000000" &
		"011001110100000001" &
		"00000000000000000000" &
		"011000110010000001" &
		"00000000000000000000" &
		"1111110000001001" &
		"00000000000000000000" &
		"01111010101111110" &
		"00000000000000000000" &
		"0110010011100000" &
		"00000000000000000000" &
		"011100110111010001" &
		"00000000000000000000" &
		"011101000111100011" &
		"00000000000000000000" &
		"11111111011001011" &
		"00000000000000000000" &
		"001101010101111001" &
		"00000000000000000000" &
		"0111111011000110" &
		"00000000000000000000" &
		"00101001100000011" &
		"00000000000000000000" &
		"0011000101110100" &
		"00000000000000000000" &
		"001111110100010101" &
		"00000000000000000000" &
		"0010010011100011" &
		"00000000000000000000" &
		"111101011101000011" &
		"00000000000000000000" &
		"00110110011" &
		"00000000000000000000" &
		"101011001011110000" &
		"00000000000000000000" &
		"1011111100001010" &
		"00000000000000000000" &
		"01110010000100001" &
		"00000000000000000000" &
		"011010011100001011" &
		"00000000000000000000" &
		"10101100111110101" &
		"00000000000000000000" &
		"10110111101101101" &
		"00000000000000000000" &
		"011111010010010010" &
		"00000000000000000000" &
		"01110001000000" &
		"00000000000000000000" &
		"1010000110000" &
		"00000000000000000000" &
		"10100101001101001" &
		"00000000000000000000" &
		"111111101101101000" &
		"00000000000000000000" &
		"011010001101111110" &
		"00000000000000000000" &
		"00101001010010001" &
		"00000000000000000000" &
		"111000110001101101" &
		"00000000000000000000" &
		"10111011001001100" &
		"00000000000000000000" &
		"0110110100101" &
		"00000000000000000000" &
		"00101111011010001" &
		"00000000000000000000" &
		"101001101011001001" &
		"00000000000000000000" &
		"001010101111011" &
		"00000000000000000000" &
		"00111100110000010" &
		"00000000000000000000" &
		"111000000111100011" &
		"00000000000000000000" &
		"001010110001111010" &
		"00000000000000000000" &
		"111101100000111" &
		"00000000000000000000" &
		"11111110011101110" &
		"00000000000000000000" &
		"111101010011010110" &
		"00000000000000000000" &
		"10100110100000" &
		"00000000000000000000" &
		"10100111100110011" &
		"00000000000000000000" &
		"011000010010000000" &
		"00000000000000000000" &
		"011001000010110101" &
		"00000000000000000000" &
		"111101000011011101" &
		"00000000000000000000" &
		"111000110011110001" &
		"00000000000000000000" &
		"101100010100010000" &
		"00000000000000000000" &
		"011001010011110101" &
		"00000000000000000000" &
		"001101001110100" &
		"00000000000000000000" &
		"00110100100001000" &
		"00000000000000000000" &
		"1011000000111111" &
		"00000000000000000000" &
		"111111010110110100" &
		"00000000000000000000" &
		"101111010110001000" &
		"00000000000000000000" &
		"0110111000001111" &
		"00000000000000000000" &
		"001011111011" &
		"00000000000000000000" &
		"001001011001011001" &
		"00000000000000000000" &
		"0010001011100110" &
		"00000000000000000000" &
		"101100011110001100" &
		"00000000000000000000" &
		"001001001100110110" &
		"00000000000000000000" &
		"1110000100111101" &
		"00000000000000000000" &
		"1111001101101101" &
		"00000000000000000000" &
		"011101000110111010" &
		"00000000000000000000" &
		"111000110000110011" &
		"00000000000000000000" &
		"01100110111000111" &
		"00000000000000000000" &
		"00100111101000100" &
		"00000000000000000000" &
		"00110111111100000" &
		"00000000000000000000" &
		"0010110100010001" &
		"00000000000000000000" &
		"001010110100000011" &
		"00000000000000000000" &
		"001011001111001111" &
		"00000000000000000000" &
		"01100011000111101" &
		"00000000000000000000" &
		"111001001000011001" &
		"00000000000000000000" &
		"10111011011110111" &
		"00000000000000000000" &
		"10100110111111010" &
		"00000000000000000000" &
		"101001000010011110" &
		"00000000000000000000" &
		"01100100111100101" &
		"00000000000000000000" &
		"011001101011010000" &
		"00000000000000000000" &
		"111000110101001100" &
		"00000000000000000000" &
		"10111001100011011" &
		"00000000000000000000" &
		"11100100111001001" &
		"00000000000000000000" &
		"11101000110101110" &
		"00000000000000000000" &
		"01100011100000011" &
		"00000000000000000000" &
		"1011010001101011" &
		"00000000000000000000" &
		"00101000100100000" &
		"00000000000000000000" &
		"011101101111100000" &
		"00000000000000000000" &
		"111000100101011010" &
		"00000000000000000000" &
		"101011101010001100" &
		"00000000000000000000" &
		"111111010010101011" &
		"00000000000000000000" &
		"0111101010010010" &
		"00000000000000000000" &
		"001110011000000" &
		"00000000000000000000" &
		"101110000111001000" &
		"00000000000000000000" &
		"11100101000110010" &
		"00000000000000000000" &
		"10110111110001001" &
		"00000000000000000000" &
		"001011000101000" &
		"00000000000000000000" &
		"101010000000001" &
		"00000000000000000000" &
		"0110110011000111" &
		"00000000000000000000" &
		"011001101010100" &
		"00000000000000000000" &
		"111100110110001101" &
		"00000000000000000000" &
		"01101100010110000" &
		"00000000000000000000" &
		"1110101101001111" &
		"00000000000000000000" &
		"001100010100110001" &
		"00000000000000000000" &
		"011000110111011" &
		"00000000000000000000" &
		"1010101000010111" &
		"00000000000000000000" &
		"001110100110010010" &
		"00000000000000000000" &
		"01101011101111" &
		"00000000000000000000" &
		"101100110011001000" &
		"00000000000000000000" &
		"00110101101110110" &
		"00000000000000000000" &
		"11110000000001010" &
		"00000000000000000000" &
		"011000000000110" &
		"00000000000000000000" &
		"101010100" &
		"00000000000000000000" &
		"11101101010111101" &
		"00000000000000000000" &
		"111011100001001100" &
		"00000000000000000000" &
		"111001101110011010" &
		"00000000000000000000" &
		"11111011011001111" &
		"00000000000000000000" &
		"101101000101010" &
		"00000000000000000000" &
		"101100110000000000" &
		"00000000000000000000" &
		"1110110011011111" &
		"00000000000000000000" &
		"011010001111010010" &
		"00000000000000000000" &
		"111001001101000001" &
		"00000000000000000000" &
		"001010100011101000" &
		"00000000000000000000" &
		"01101110100100001" &
		"00000000000000000000" &
		"001010110110000111" &
		"00000000000000000000" &
		"011100011011011000" &
		"00000000000000000000" &
		"101011101101100011" &
		"00000000000000000000" &
		"101011010010101100" &
		"00000000000000000000" &
		"111100010111101010" &
		"00000000000000000000" &
		"001110001010011100" &
		"00000000000000000000" &
		"11100100011101011" &
		"00000000000000000000" &
		"101011110001100000" &
		"00000000000000000000" &
		"0110011011110110" &
		"00000000000000000000" &
		"11100110000110" &
		"00000000000000000000" &
		"1111000101011" &
		"00000000000000000000" &
		"00101111001101101" &
		"00000000000000000000" &
		"101000001111001011" &
		"00000000000000000000" &
		"01100011100000001" &
		"00000000000000000000" &
		"1011100111100101" &
		"00000000000000000000" &
		"10101111001010010" &
		"00000000000000000000" &
		"01100100100000100" &
		"00000000000000000000" &
		"0010010001000111" &
		"00000000000000000000" &
		"111000101111100" &
		"00000000000000000000" &
		"001110101111100100" &
		"00000000000000000000" &
		"101111011001010000" &
		"00000000000000000000" &
		"011011011000001101" &
		"00000000000000000000" &
		"1010110110111" &
		"00000000000000000000" &
		"01100000001101100" &
		"00000000000000000000" &
		"001101010000001001" &
		"00000000000000000000" &
		"01111111010100000" &
		"00000000000000000000" &
		"11110101010011011" &
		"00000000000000000000" &
		"111010001010001111" &
		"00000000000000000000" &
		"011010000110" &
		"00000000000000000000" &
		"11101001011110000" &
		"00000000000000000000" &
		"01110100110101111" &
		"00000000000000000000" &
		"011101111010011110" &
		"00000000000000000000" &
		"1111111100000100" &
		"00000000000000000000" &
		"1111110111001100" &
		"00000000000000000000" &
		"001011111110110" &
		"00000000000000000000" &
		"10110011101001111" &
		"00000000000000000000" &
		"10110011110111101" &
		"00000000000000000000" &
		"0110101011001101" &
		"00000000000000000000" &
		"101010001101110111" &
		"00000000000000000000" &
		"011010110000110100" &
		"00000000000000000000" &
		"10110111000110001" &
		"00000000000000000000" &
		"11101000000001000" &
		"00000000000000000000" &
		"1111100111001100" &
		"00000000000000000000" &
		"11111011011001000" &
		"00000000000000000000" &
		"001011010111011111" &
		"00000000000000000000" &
		"001111001100000" &
		"00000000000000000000" &
		"001111011001001101" &
		"00000000000000000000" &
		"001010100010000011" &
		"00000000000000000000" &
		"01110111010110111" &
		"00000000000000000000" &
		"001000101010010000" &
		"00000000000000000000" &
		"0011101110001010" &
		"00000000000000000000" &
		"011110001101111111" &
		"00000000000000000000" &
		"01110011101101" &
		"00000000000000000000" &
		"01101000001111110" &
		"00000000000000000000" &
		"0010101001010110" &
		"00000000000000000000" &
		"00111101001100100" &
		"00000000000000000000" &
		"00101010111110010" &
		"00000000000000000000" &
		"11101000101010000" &
		"00000000000000000000" &
		"00110001000000101" &
		"00000000000000000000" &
		"10110000110111010" &
		"00000000000000000000" &
		"101110011110101011" &
		"00000000000000000000" &
		"1011001101101010" &
		"00000000000000000000" &
		"011010101111010010" &
		"00000000000000000000" &
		"1110110011000011" &
		"00000000000000000000" &
		"001111001010001001" &
		"00000000000000000000" &
		"011101000010100110" &
		"00000000000000000000" &
		"1011110011100011" &
		"00000000000000000000" &
		"11101101000000011" &
		"00000000000000000000" &
		"10101111011110110" &
		"00000000000000000000" &
		"0011101010111011" &
		"00000000000000000000" &
		"11111000000001100" &
		"00000000000000000000" &
		"101110011010110010" &
		"00000000000000000000" &
		"001000011010000100" &
		"00000000000000000000" &
		"101110011111100011" &
		"00000000000000000000" &
		"001010100100000101" &
		"00000000000000000000" &
		"011110100010111110" &
		"00000000000000000000" &
		"00100110011100011" &
		"00000000000000000000" &
		"111000001110110111" &
		"00000000000000000000" &
		"01100001110100111" &
		"00000000000000000000" &
		"10101110011100" &
		"00000000000000000000" &
		"111010001100111000" &
		"00000000000000000000" &
		"00100000110110001" &
		"00000000000000000000" &
		"00101110000010111" &
		"00000000000000000000" &
		"1111101100000100" &
		"00000000000000000000" &
		"11100110110101001" &
		"00000000000000000000" &
		"01101100000110" &
		"00000000000000000000" &
		"0010110110001101" &
		"00000000000000000000" &
		"10101001100000101" &
		"00000000000000000000" &
		"111001100101001110" &
		"00000000000000000000" &
		"10100000111101101" &
		"00000000000000000000" &
		"00111100011000011" &
		"00000000000000000000" &
		"001111100111110010" &
		"00000000000000000000" &
		"0111110010111110" &
		"00000000000000000000" &
		"1110011101011001" &
		"00000000000000000000" &
		"011010101111010101" &
		"00000000000000000000" &
		"011101000001010100" &
		"00000000000000000000" &
		"01111010010010101" &
		"00000000000000000000" &
		"011111100101011000" &
		"00000000000000000000" &
		"001111011010111010" &
		"00000000000000000000" &
		"1110000101100100" &
		"00000000000000000000" &
		"001011011111110010" &
		"00000000000000000000" &
		"0110001011101101" &
		"00000000000000000000" &
		"1110010100010100" &
		"00000000000000000000" &
		"111101000111000001" &
		"00000000000000000000" &
		"1111011001111010" &
		"00000000000000000000" &
		"11100001001001001" &
		"00000000000000000000" &
		"111111010011001001" &
		"00000000000000000000" &
		"11100011000010110" &
		"00000000000000000000" &
		"00101011011100111" &
		"00000000000000000000" &
		"11101001110010110" &
		"00000000000000000000" &
		"001000101010111100" &
		"00000000000000000000" &
		"111011001001000000" &
		"00000000000000000000" &
		"00101000110011000" &
		"00000000000000000000" &
		"101001000000101101" &
		"00000000000000000000" &
		"111000010100111111" &
		"00000000000000000000" &
		"10110101001100001" &
		"00000000000000000000" &
		"00111011001001001" &
		"00000000000000000000" &
		"101001100110001011" &
		"00000000000000000000" &
		"001001011010" &
		"00000000000000000000" &
		"10101111001111" &
		"00000000000000000000" &
		"001001010011001001" &
		"00000000000000000000" &
		"1010100001101101" &
		"00000000000000000000" &
		"0110111000000001" &
		"00000000000000000000" &
		"111100111010001111" &
		"00000000000000000000" &
		"0110010101110100" &
		"00000000000000000000" &
		"01100000010111100" &
		"00000000000000000000" &
		"10100000100100011" &
		"00000000000000000000" &
		"11111111111101100" &
		"00000000000000000000" &
		"011001010100010101" &
		"00000000000000000000" &
		"1010100100111" &
		"00000000000000000000" &
		"001101101100" &
		"00000000000000000000" &
		"10101010101110" &
		"00000000000000000000" &
		"101111011100010" &
		"00000000000000000000" &
		"101110100001011000" &
		"00000000000000000000" &
		"00110111110011110" &
		"00000000000000000000" &
		"101000110101101110" &
		"00000000000000000000" &
		"001111101011011011" &
		"00000000000000000000" &
		"101011100110001111" &
		"00000000000000000000" &
		"1010001101100010" &
		"00000000000000000000" &
		"011100101011100011" &
		"00000000000000000000" &
		"01110101000110000" &
		"00000000000000000000" &
		"001111101001000000" &
		"00000000000000000000" &
		"011111101101010111" &
		"00000000000000000000" &
		"011000111111101000" &
		"00000000000000000000" &
		"111000010110010" &
		"00000000000000000000" &
		"0011001111111001" &
		"00000000000000000000" &
		"11110001011000100" &
		"00000000000000000000" &
		"001101110001000101" &
		"00000000000000000000" &
		"00111111001110111" &
		"00000000000000000000" &
		"10101101001100111" &
		"00000000000000000000" &
		"00110111000101001" &
		"00000000000000000000" &
		"0111110001111000" &
		"00000000000000000000" &
		"101110100101000001" &
		"00000000000000000000" &
		"011011010111000000" &
		"00000000000000000000" &
		"101110100111111010" &
		"00000000000000000000" &
		"0011101100001" &
		"00000000000000000000" &
		"10101001101000101" &
		"00000000000000000000" &
		"001011110010001000" &
		"00000000000000000000" &
		"101010110000010101" &
		"00000000000000000000" &
		"00110000110001" &
		"00000000000000000000" &
		"11111000101100001" &
		"00000000000000000000" &
		"00100110000110111" &
		"00000000000000000000" &
		"111111010010011110" &
		"00000000000000000000" &
		"001000101101110110" &
		"00000000000000000000" &
		"111001101101100111" &
		"00000000000000000000" &
		"001011011111101000" &
		"00000000000000000000" &
		"001110111101001010" &
		"00000000000000000000" &
		"111010010110011100" &
		"00000000000000000000" &
		"0110010000010" &
		"00000000000000000000" &
		"101101010000101011" &
		"00000000000000000000" &
		"11110000010100011" &
		"00000000000000000000" &
		"01101111111101101" &
		"00000000000000000000" &
		"1011101111011110" &
		"00000000000000000000" &
		"00111011110111001" &
		"00000000000000000000" &
		"011111000101100000" &
		"00000000000000000000" &
		"1111000010111010" &
		"00000000000000000000" &
		"10111011100001000" &
		"00000000000000000000" &
		"11110000111000000" &
		"00000000000000000000" &
		"111111001110001011" &
		"00000000000000000000" &
		"1010001100010" &
		"00000000000000000000" &
		"111100110111111000" &
		"00000000000000000000" &
		"1111110011001" &
		"00000000000000000000" &
		"001000010101100000" &
		"00000000000000000000" &
		"00110100011010101" &
		"00000000000000000000" &
		"101101000111000111" &
		"00000000000000000000" &
		"011101100000100111" &
		"00000000000000000000" &
		"1010100100" &
		"00000000000000000000" &
		"001010000110000011" &
		"00000000000000000000" &
		"001100000010110010" &
		"00000000000000000000" &
		"01100010101" &
		"00000000000000000000" &
		"001101001010010" &
		"00000000000000000000" &
		"101000111010101001" &
		"00000000000000000000" &
		"00110001010110010" &
		"00000000000000000000" &
		"011001101110111" &
		"00000000000000000000" &
		"001011110001110100" &
		"00000000000000000000" &
		"111101010111001011" &
		"00000000000000000000" &
		"11111011111101111" &
		"00000000000000000000" &
		"01100101000101110" &
		"00000000000000000000" &
		"001001001101101100" &
		"00000000000000000000" &
		"011010001010000000" &
		"00000000000000000000" &
		"011110011000110100" &
		"00000000000000000000" &
		"00100111100011000" &
		"00000000000000000000" &
		"111011000100001100" &
		"00000000000000000000" &
		"10111010110010101" &
		"00000000000000000000" &
		"0111011011100010" &
		"00000000000000000000" &
		"10101000011100001" &
		"00000000000000000000" &
		"111100001010110100" &
		"00000000000000000000" &
		"111000111001011001" &
		"00000000000000000000" &
		"101011010011101010" &
		"00000000000000000000" &
		"011101100101100010" &
		"00000000000000000000" &
		"011111110010000001" &
		"00000000000000000000" &
		"001000100000000010" &
		"00000000000000000000" &
		"00111111111" &
		"00000000000000000000" &
		"01111110101110110" &
		"00000000000000000000" &
		"101100011100111010" &
		"00000000000000000000" &
		"11100110101000100" &
		"00000000000000000000" &
		"1111010111001010" &
		"00000000000000000000" &
		"1111110010010010" &
		"00000000000000000000" &
		"011111011001011111" &
		"00000000000000000000" &
		"101010110000" &
		"00000000000000000000" &
		"01101101001100001" &
		"00000000000000000000" &
		"011101011011011110" &
		"00000000000000000000" &
		"0111111110000000" &
		"00000000000000000000" &
		"011010100110111011" &
		"00000000000000000000" &
		"011011000101011000" &
		"00000000000000000000" &
		"111000001101101" &
		"00000000000000000000" &
		"001101000000001111" &
		"00000000000000000000" &
		"011111010110010111" &
		"00000000000000000000" &
		"1110000101111" &
		"00000000000000000000" &
		"011111011101110011" &
		"00000000000000000000" &
		"001010010000001010" &
		"00000000000000000000" &
		"101011100111010" &
		"00000000000000000000" &
		"00101001101100" &
		"00000000000000000000" &
		"111010001101000100" &
		"00000000000000000000" &
		"101101100111101110" &
		"00000000000000000000" &
		"101111010110101111" &
		"00000000000000000000" &
		"011011010011110111" &
		"00000000000000000000" &
		"00110000101101000" &
		"00000000000000000000" &
		"101011111100011001" &
		"00000000000000000000" &
		"111011011111001" &
		"00000000000000000000" &
		"111001011110100001" &
		"00000000000000000000" &
		"101101001010011101" &
		"00000000000000000000" &
		"001110111100010" &
		"00000000000000000000" &
		"1110010111001010" &
		"00000000000000000000" &
		"101001111000000" &
		"00000000000000000000" &
		"01101101100101000" &
		"00000000000000000000" &
		"011100110111001111" &
		"00000000000000000000" &
		"101101010000000101" &
		"00000000000000000000" &
		"1011111101010000" &
		"00000000000000000000" &
		"101100000010110" &
		"00000000000000000000" &
		"11101111010100001" &
		"00000000000000000000" &
		"111101010001101101" &
		"00000000000000000000" &
		"01101111000111010" &
		"00000000000000000000" &
		"011011101110111010" &
		"00000000000000000000" &
		"0010100010000001" &
		"00000000000000000000" &
		"001001001110011001" &
		"00000000000000000000" &
		"001110100101100100" &
		"00000000000000000000" &
		"0110110110001100" &
		"00000000000000000000" &
		"11100010010111111" &
		"00000000000000000000" &
		"0010111111110001" &
		"00000000000000000000" &
		"101001100010000010" &
		"00000000000000000000" &
		"00110110110010001" &
		"00000000000000000000" &
		"01100111100110110" &
		"00000000000000000000" &
		"101000111101100100" &
		"00000000000000000000" &
		"111010101001010101" &
		"00000000000000000000" &
		"1111011111101101" &
		"00000000000000000000" &
		"001001011101011" &
		"00000000000000000000" &
		"001001110001101000" &
		"00000000000000000000" &
		"011110111100011111" &
		"00000000000000000000" &
		"101111010010100110" &
		"00000000000000000000" &
		"011101010101010101" &
		"00000000000000000000" &
		"10101010110101100" &
		"00000000000000000000" &
		"101100100011010001" &
		"00000000000000000000" &
		"111000110100010100" &
		"00000000000000000000" &
		"00101110001010100" &
		"00000000000000000000" &
		"11110010111000" &
		"00000000000000000000" &
		"00111110111001100" &
		"00000000000000000000" &
		"111111101101000001" &
		"00000000000000000000" &
		"10110010110000000" &
		"00000000000000000000" &
		"00111010010010010" &
		"00000000000000000000" &
		"111110010000100111" &
		"00000000000000000000" &
		"101111100010101011" &
		"00000000000000000000" &
		"0011100110100" &
		"00000000000000000000" &
		"011011110110111101" &
		"00000000000000000000" &
		"01100010001011111" &
		"00000000000000000000" &
		"11101001111001001" &
		"00000000000000000000" &
		"111010011001101101" &
		"00000000000000000000" &
		"001010101000011111" &
		"00000000000000000000" &
		"101111100101000111" &
		"00000000000000000000" &
		"101010100001101100" &
		"00000000000000000000" &
		"011110001110100111" &
		"00000000000000000000" &
		"011001000110100001" &
		"00000000000000000000" &
		"111101001110011101" &
		"00000000000000000000" &
		"101010001100111011" &
		"00000000000000000000" &
		"01111100000100011" &
		"00000000000000000000" &
		"001111010100100010" &
		"00000000000000000000" &
		"001101100000001001" &
		"00000000000000000000" &
		"0010100000010100" &
		"00000000000000000000" &
		"001010101111001100" &
		"00000000000000000000" &
		"011000101001011001" &
		"00000000000000000000" &
		"0011100101" &
		"00000000000000000000" &
		"001100010100000101" &
		"00000000000000000000" &
		"11110110011101110" &
		"00000000000000000000" &
		"101011110100001" &
		"00000000000000000000" &
		"111001100011110101" &
		"00000000000000000000" &
		"1111111110000000" &
		"00000000000000000000" &
		"111000100010111" &
		"00000000000000000000" &
		"00111101100010001" &
		"00000000000000000000" &
		"10111000110011001" &
		"00000000000000000000" &
		"1111010001011000" &
		"00000000000000000000" &
		"1111111011010000" &
		"00000000000000000000" &
		"101101011110100101" &
		"00000000000000000000" &
		"111101100000001101" &
		"00000000000000000000" &
		"111100000011000" &
		"00000000000000000000" &
		"001100111110010100" &
		"00000000000000000000" &
		"111000011100010011" &
		"00000000000000000000" &
		"00100101111010011" &
		"00000000000000000000" &
		"001000010010110001" &
		"00000000000000000000" &
		"11101001110110110" &
		"00000000000000000000" &
		"01101100101101000" &
		"00000000000000000000" &
		"001001010100010101" &
		"00000000000000000000" &
		"001011111101101011" &
		"00000000000000000000" &
		"001000011100000001" &
		"00000000000000000000" &
		"011001011110110000" &
		"00000000000000000000" &
		"001100000110100" &
		"00000000000000000000" &
		"101101111011111" &
		"00000000000000000000" &
		"1011000111000010" &
		"00000000000000000000" &
		"1010001011000" &
		"00000000000000000000" &
		"01110110100101001" &
		"00000000000000000000" &
		"10110111001101110" &
		"00000000000000000000" &
		"01101011001101011" &
		"00000000000000000000" &
		"0011001011010" &
		"00000000000000000000" &
		"011011010101111001" &
		"00000000000000000000" &
		"111011101101110001" &
		"00000000000000000000" &
		"001101011010110111" &
		"00000000000000000000" &
		"111111000110110" &
		"00000000000000000000" &
		"101111001001101110" &
		"00000000000000000000" &
		"0110000001111011" &
		"00000000000000000000" &
		"001010111111100100" &
		"00000000000000000000" &
		"111100000100001110" &
		"00000000000000000000" &
		"001110010110010010" &
		"00000000000000000000" &
		"011100101101110100" &
		"00000000000000000000" &
		"111010010011101000" &
		"00000000000000000000" &
		"01111000010001" &
		"00000000000000000000" &
		"01101110010101100" &
		"00000000000000000000" &
		"111001101011110111" &
		"00000000000000000000" &
		"111100011101110001" &
		"00000000000000000000" &
		"0011011001110000" &
		"00000000000000000000" &
		"011110001011101011" &
		"00000000000000000000" &
		"01111001101110111" &
		"00000000000000000000" &
		"0011100011101011" &
		"00000000000000000000" &
		"11101010011100111" &
		"00000000000000000000" &
		"101110001101100010" &
		"00000000000000000000" &
		"10111010010100001" &
		"00000000000000000000" &
		"0110111010100010" &
		"00000000000000000000" &
		"01110110101100011" &
		"00000000000000000000" &
		"1111101000100011" &
		"00000000000000000000" &
		"011010001101110000" &
		"00000000000000000000" &
		"0010011100100001" &
		"00000000000000000000" &
		"111010010010000010" &
		"00000000000000000000" &
		"0110110001101110" &
		"00000000000000000000" &
		"101000101111111110" &
		"00000000000000000000" &
		"11101010111100111" &
		"00000000000000000000" &
		"00100011000110" &
		"00000000000000000000" &
		"011010011001100000" &
		"00000000000000000000" &
		"00110011010011100" &
		"00000000000000000000" &
		"001011010011100001" &
		"00000000000000000000" &
		"10100100101110011" &
		"00000000000000000000" &
		"0111100111001101" &
		"00000000000000000000" &
		"111101011011111111" &
		"00000000000000000000" &
		"10110001010001101" &
		"00000000000000000000" &
		"00100001011010" &
		"00000000000000000000" &
		"0011011110101101" &
		"00000000000000000000" &
		"101011001101101101" &
		"00000000000000000000" &
		"11100100101010110" &
		"00000000000000000000" &
		"001110000001010000" &
		"00000000000000000000" &
		"101100001001011010" &
		"00000000000000000000" &
		"101100100100000100" &
		"00000000000000000000" &
		"111000010100100010" &
		"00000000000000000000" &
		"1010000100101011" &
		"00000000000000000000" &
		"101111001100001000" &
		"00000000000000000000" &
		"111101000000100000" &
		"00000000000000000000" &
		"01100100000000110" &
		"00000000000000000000" &
		"011100010100000001" &
		"00000000000000000000" &
		"011011110110011000" &
		"00000000000000000000" &
		"111100100110101000" &
		"00000000000000000000" &
		"001110111111011010" &
		"00000000000000000000" &
		"001010001110010001" &
		"00000000000000000000" &
		"001000010011110010" &
		"00000000000000000000" &
		"101001111000111010" &
		"00000000000000000000" &
		"1010010101011010" &
		"00000000000000000000" &
		"0010101010010100" &
		"00000000000000000000" &
		"001100111101101010" &
		"00000000000000000000" &
		"101011100011010" &
		"00000000000000000000" &
		"011111011000100110" &
		"00000000000000000000" &
		"001110100101111000" &
		"00000000000000000000" &
		"00101101001100000" &
		"00000000000000000000" &
		"001010011111111011" &
		"00000000000000000000" &
		"10110100010001101" &
		"00000000000000000000" &
		"001011111100101010" &
		"00000000000000000000" &
		"10110101011000000" &
		"00000000000000000000" &
		"0011101001111010" &
		"00000000000000000000" &
		"101100111100" &
		"00000000000000000000" &
		"0111000000100010" &
		"00000000000000000000" &
		"1011010011001010" &
		"00000000000000000000" &
		"011010111111100101" &
		"00000000000000000000" &
		"01110001100011011" &
		"00000000000000000000" &
		"011100011001100" &
		"00000000000000000000" &
		"011100000111101" &
		"00000000000000000000" &
		"011010001110000100" &
		"00000000000000000000" &
		"0011111111100000" &
		"00000000000000000000" &
		"00101000101111101" &
		"00000000000000000000" &
		"111111110010101110" &
		"00000000000000000000" &
		"101010101010101000" &
		"00000000000000000000" &
		"011110100110000101" &
		"00000000000000000000" &
		"001010101100110101" &
		"00000000000000000000" &
		"10101100000101100" &
		"00000000000000000000" &
		"11110101011110111" &
		"00000000000000000000" &
		"001111100101000101" &
		"00000000000000000000" &
		"101011111000100011" &
		"00000000000000000000" &
		"1110110010000011" &
		"00000000000000000000" &
		"101000011111110010" &
		"00000000000000000000" &
		"011010100010011" &
		"00000000000000000000" &
		"101010101110010001" &
		"00000000000000000000" &
		"011111100010100" &
		"00000000000000000000" &
		"101001101110101100" &
		"00000000000000000000" &
		"101111000010100100" &
		"00000000000000000000" &
		"101010010001010001" &
		"00000000000000000000" &
		"101010100010101101" &
		"00000000000000000000" &
		"01101101001011001" &
		"00000000000000000000" &
		"11100000010000100" &
		"00000000000000000000" &
		"1011011101011" &
		"00000000000000000000" &
		"001111110101010110" &
		"00000000000000000000" &
		"001001100101010000" &
		"00000000000000000000" &
		"001111111001" &
		"00000000000000000000" &
		"111001010101000011" &
		"00000000000000000000" &
		"00110100111111101" &
		"00000000000000000000" &
		"11111010000110011" &
		"00000000000000000000" &
		"1111110101011" &
		"00000000000000000000" &
		"011101110101000011" &
		"00000000000000000000" &
		"10111100001110001" &
		"00000000000000000000" &
		"011101100000010101" &
		"00000000000000000000" &
		"0010001001111100" &
		"00000000000000000000" &
		"001101011001001100" &
		"00000000000000000000" &
		"0011100100100000" &
		"00000000000000000000" &
		"11111010000011010" &
		"00000000000000000000" &
		"1111110011101100" &
		"00000000000000000000" &
		"11110111010" &
		"00000000000000000000" &
		"111001111010001011" &
		"00000000000000000000" &
		"011000110100110111" &
		"00000000000000000000" &
		"001111001100100001" &
		"00000000000000000000" &
		"10111000011111110" &
		"00000000000000000000" &
		"011011001111010010" &
		"00000000000000000000" &
		"011101000110110" &
		"00000000000000000000" &
		"111000001111100010" &
		"00000000000000000000" &
		"10111100010001110" &
		"00000000000000000000" &
		"011110101100011000" &
		"00000000000000000000" &
		"111001001010100111" &
		"00000000000000000000" &
		"111000111011101111" &
		"00000000000000000000" &
		"1111010110111100" &
		"00000000000000000000" &
		"1011100111000101" &
		"00000000000000000000" &
		"0111001000110110" &
		"00000000000000000000" &
		"00111000011101110" &
		"00000000000000000000" &
		"111011111001100" &
		"00000000000000000000" &
		"011100110100100001" &
		"00000000000000000000" &
		"011111010100111000" &
		"00000000000000000000" &
		"001001001101011111" &
		"00000000000000000000" &
		"001111110011000010" &
		"00000000000000000000" &
		"101100001010111000" &
		"00000000000000000000" &
		"001001000101111010" &
		"00000000000000000000" &
		"0111100101000010" &
		"00000000000000000000" &
		"001110101110110001" &
		"00000000000000000000" &
		"111101111100000110" &
		"00000000000000000000" &
		"011001100001010111" &
		"00000000000000000000" &
		"111000011100111101" &
		"00000000000000000000" &
		"11101010101110111" &
		"00000000000000000000" &
		"011011101001011000" &
		"00000000000000000000" &
		"11110111100111001" &
		"00000000000000000000" &
		"111101010011101000" &
		"00000000000000000000" &
		"001100010110010101" &
		"00000000000000000000" &
		"011011101100101110" &
		"00000000000000000000" &
		"111000000100011010" &
		"00000000000000000000" &
		"10111000110001011" &
		"00000000000000000000" &
		"111111000111" &
		"00000000000000000000" &
		"101010001001010010" &
		"00000000000000000000" &
		"101001010101111111" &
		"00000000000000000000" &
		"011111010110000100" &
		"00000000000000000000" &
		"11100111000110110" &
		"00000000000000000000" &
		"111111001001011001" &
		"00000000000000000000" &
		"111001100001001101" &
		"00000000000000000000" &
		"111000010100100000" &
		"00000000000000000000" &
		"1010011110010101" &
		"00000000000000000000" &
		"001011000100110100" &
		"00000000000000000000" &
		"001101100000010010" &
		"00000000000000000000" &
		"111101010100110010" &
		"00000000000000000000" &
		"01111010110010" &
		"00000000000000000000" &
		"1110000011001111" &
		"00000000000000000000" &
		"1111001110001000" &
		"00000000000000000000" &
		"1011011000101" &
		"00000000000000000000" &
		"1011010101000010" &
		"00000000000000000000" &
		"111001111000000101" &
		"00000000000000000000" &
		"101000110110100010" &
		"00000000000000000000" &
		"0110011010000101" &
		"00000000000000000000" &
		"101000001010111111" &
		"00000000000000000000" &
		"001110101001010111" &
		"00000000000000000000" &
		"11101111010111111" &
		"00000000000000000000" &
		"101101100001110001" &
		"00000000000000000000" &
		"111100110100100111" &
		"00000000000000000000" &
		"1111010101110001" &
		"00000000000000000000" &
		"1010001111011011" &
		"00000000000000000000" &
		"011000000011010101" &
		"00000000000000000000" &
		"101001010000000010" &
		"00000000000000000000" &
		"0010110000010000" &
		"00000000000000000000" &
		"00111101011101101" &
		"00000000000000000000" &
		"01110000110011000" &
		"00000000000000000000" &
		"11101111010100111" &
		"00000000000000000000" &
		"0110110111111100" &
		"00000000000000000000" &
		"101101010001111011" &
		"00000000000000000000" &
		"00100100100011110" &
		"00000000000000000000" &
		"01100011111001111" &
		"00000000000000000000" &
		"001010000101010011" &
		"00000000000000000000" &
		"101000001010101011" &
		"00000000000000000000" &
		"011011111100111110" &
		"00000000000000000000" &
		"101010101011101" &
		"00000000000000000000" &
		"011010101111110100" &
		"00000000000000000000" &
		"01101101000101101" &
		"00000000000000000000" &
		"00100000011011110" &
		"00000000000000000000" &
		"011110001101101000" &
		"00000000000000000000" &
		"111101110111000000" &
		"00000000000000000000" &
		"11101000111110101" &
		"00000000000000000000" &
		"001010000010011010" &
		"00000000000000000000" &
		"101101000101010111" &
		"00000000000000000000" &
		"1010001100111110" &
		"00000000000000000000" &
		"001101100001100" &
		"00000000000000000000" &
		"101011000100101110" &
		"00000000000000000000" &
		"11100011010010101" &
		"00000000000000000000" &
		"101110001111111010" &
		"00000000000000000000" &
		"1010100000101001" &
		"00000000000000000000" &
		"01101111111110010" &
		"00000000000000000000" &
		"01110010100011100" &
		"00000000000000000000" &
		"10100001111111110" &
		"00000000000000000000" &
		"101100111010010001" &
		"00000000000000000000" &
		"001101111111101001" &
		"00000000000000000000" &
		"0110101101010101" &
		"00000000000000000000" &
		"001100110101011001" &
		"00000000000000000000" &
		"011100011000110011" &
		"00000000000000000000" &
		"111001001111001100" &
		"00000000000000000000" &
		"1010011111011010" &
		"00000000000000000000" &
		"011100100111011100" &
		"00000000000000000000" &
		"001011111010100110" &
		"00000000000000000000" &
		"01110100010001100" &
		"00000000000000000000" &
		"011010011001101101" &
		"00000000000000000000" &
		"111110000000011110" &
		"00000000000000000000" &
		"011001110010111001" &
		"00000000000000000000" &
		"001001101011101110" &
		"00000000000000000000" &
		"011011110001001110" &
		"00000000000000000000" &
		"001101101001010010" &
		"00000000000000000000" &
		"111000111101100110" &
		"00000000000000000000" &
		"111101010000000001" &
		"00000000000000000000" &
		"101000000010101110" &
		"00000000000000000000" &
		"001000100011000111" &
		"00000000000000000000" &
		"111010000000000100" &
		"00000000000000000000" &
		"111010100010111010" &
		"00000000000000000000" &
		"00101010001000000" &
		"00000000000000000000" &
		"111110111101010000" &
		"00000000000000000000" &
		"0110000111011010" &
		"00000000000000000000" &
		"0011010000011001" &
		"00000000000000000000" &
		"11101101101010010" &
		"00000000000000000000" &
		"00100100100111" &
		"00000000000000000000" &
		"101001101100111110" &
		"00000000000000000000" &
		"111010010010001000" &
		"00000000000000000000" &
		"0010000110111001" &
		"00000000000000000000" &
		"011010001110011110" &
		"00000000000000000000" &
		"011010101010001010" &
		"00000000000000000000" &
		"001011000100000" &
		"00000000000000000000" &
		"11101001000110011" &
		"00000000000000000000" &
		"10110011101101" &
		"00000000000000000000" &
		"101000011000111100" &
		"00000000000000000000" &
		"011100100011110111" &
		"00000000000000000000" &
		"1110100010001110" &
		"00000000000000000000" &
		"01101011011010" &
		"00000000000000000000" &
		"111010110101100010" &
		"00000000000000000000" &
		"10101101011001100" &
		"00000000000000000000" &
		"111001001110011111" &
		"00000000000000000000" &
		"111101001101100010" &
		"00000000000000000000" &
		"111011101001111111" &
		"00000000000000000000" &
		"10110011101011" &
		"00000000000000000000" &
		"101110000100011001" &
		"00000000000000000000" &
		"10100011001101100" &
		"00000000000000000000" &
		"111100111010111011" &
		"00000000000000000000" &
		"111111010010111010" &
		"00000000000000000000" &
		"0110010011101010" &
		"00000000000000000000" &
		"01110011110001100" &
		"00000000000000000000" &
		"001010000000110100" &
		"00000000000000000000" &
		"111011010101100111" &
		"00000000000000000000" &
		"011111010010110000" &
		"00000000000000000000" &
		"001100101111011000" &
		"00000000000000000000" &
		"10101110111100101" &
		"00000000000000000000" &
		"011010011100001000" &
		"00000000000000000000" &
		"011110110000110111" &
		"00000000000000000000" &
		"001111100001110100" &
		"00000000000000000000" &
		"111100101100101100" &
		"00000000000000000000" &
		"11100100111010000" &
		"00000000000000000000" &
		"101011001101101" &
		"00000000000000000000" &
		"1110100100111100" &
		"00000000000000000000" &
		"011000110001110011" &
		"00000000000000000000" &
		"101011011011110" &
		"00000000000000000000" &
		"001011110100100000" &
		"00000000000000000000" &
		"001000010111100001" &
		"00000000000000000000" &
		"001010010111110100" &
		"00000000000000000000" &
		"01111110001011000" &
		"00000000000000000000" &
		"001001011111101111" &
		"00000000000000000000" &
		"011110101101110111" &
		"00000000000000000000" &
		"101100100101110010" &
		"00000000000000000000" &
		"00100111101001" &
		"00000000000000000000" &
		"011011101011110110" &
		"00000000000000000000" &
		"00100101111111001" &
		"00000000000000000000" &
		"111100110100000" &
		"00000000000000000000" &
		"011010100001111000" &
		"00000000000000000000" &
		"10100011100" &
		"00000000000000000000" &
		"111010100010000" &
		"00000000000000000000" &
		"111100111101001011" &
		"00000000000000000000" &
		"101000010000110010" &
		"00000000000000000000" &
		"101110101110110110" &
		"00000000000000000000" &
		"11100100011011000" &
		"00000000000000000000" &
		"111000101010000111" &
		"00000000000000000000" &
		"11101000100101011" &
		"00000000000000000000" &
		"111111010010111011" &
		"00000000000000000000" &
		"001100101011101100" &
		"00000000000000000000" &
		"01100101010111001" &
		"00000000000000000000" &
		"011110111010101111" &
		"00000000000000000000" &
		"00111011001000111" &
		"00000000000000000000" &
		"111100011010001101" &
		"00000000000000000000" &
		"001101100000111101" &
		"00000000000000000000" &
		"011011011001110110" &
		"00000000000000000000" &
		"101000110110111000" &
		"00000000000000000000" &
		"1011011100011" &
		"00000000000000000000" &
		"00100011110011100" &
		"00000000000000000000" &
		"10101101110101001" &
		"00000000000000000000" &
		"00100010101010010" &
		"00000000000000000000" &
		"011110010101000001" &
		"00000000000000000000" &
		"001000100010111000" &
		"00000000000000000000" &
		"10101101100101110" &
		"00000000000000000000" &
		"101001111011010011" &
		"00000000000000000000" &
		"1010000101100010" &
		"00000000000000000000" &
		"001000011010111100" &
		"00000000000000000000" &
		"10110011110111001" &
		"00000000000000000000" &
		"101100000110110110" &
		"00000000000000000000" &
		"001011111010001111" &
		"00000000000000000000" &
		"101111001010000111" &
		"00000000000000000000" &
		"011110001110010" &
		"00000000000000000000" &
		"011111101011010110" &
		"00000000000000000000" &
		"10100001001" &
		"00000000000000000000" &
		"101110010101010000" &
		"00000000000000000000" &
		"11100001011100001" &
		"00000000000000000000" &
		"1011110110011000" &
		"00000000000000000000" &
		"00111111101000000" &
		"00000000000000000000" &
		"00100111010001111" &
		"00000000000000000000" &
		"01111000011010010" &
		"00000000000000000000" &
		"11100110011101110" &
		"00000000000000000000" &
		"011100000110111110" &
		"00000000000000000000" &
		"1010011100001110" &
		"00000000000000000000" &
		"111000011101100111" &
		"00000000000000000000" &
		"11111110010010" &
		"00000000000000000000" &
		"01101110101101101" &
		"00000000000000000000" &
		"101111001010101000" &
		"00000000000000000000" &
		"10110111100011011" &
		"00000000000000000000" &
		"001111010011100010" &
		"00000000000000000000" &
		"011001101111101100" &
		"00000000000000000000" &
		"001001001111101110" &
		"00000000000000000000" &
		"11111011110000010" &
		"00000000000000000000" &
		"101010010010011000" &
		"00000000000000000000" &
		"0010111010011001" &
		"00000000000000000000" &
		"101011001100100000" &
		"00000000000000000000" &
		"001000111111111000" &
		"00000000000000000000" &
		"00101000010100101" &
		"00000000000000000000" &
		"10110101010110000" &
		"00000000000000000000" &
		"01110000000110100" &
		"00000000000000000000" &
		"011010010001111011" &
		"00000000000000000000" &
		"001000101100011100" &
		"00000000000000000000" &
		"101100100111100101" &
		"00000000000000000000" &
		"10100101001000000" &
		"00000000000000000000" &
		"011011111100100001" &
		"00000000000000000000" &
		"111111000110000" &
		"00000000000000000000" &
		"001010011101100100" &
		"00000000000000000000" &
		"11101001110111100" &
		"00000000000000000000" &
		"111010010011111010" &
		"00000000000000000000" &
		"10110101010111" &
		"00000000000000000000" &
		"00101001000000000" &
		"00000000000000000000" &
		"11100011100101100" &
		"00000000000000000000" &
		"101110000001011101" &
		"00000000000000000000" &
		"011110010110100000" &
		"00000000000000000000" &
		"101011100100101000" &
		"00000000000000000000" &
		"0111110011101111" &
		"00000000000000000000" &
		"111110010001010010" &
		"00000000000000000000" &
		"001111101101000" &
		"00000000000000000000" &
		"0010010011100011" &
		"00000000000000000000" &
		"101111000010111100" &
		"00000000000000000000" &
		"00100111101000011" &
		"00000000000000000000" &
		"011011010010010011" &
		"00000000000000000000" &
		"0111010000110110" &
		"00000000000000000000" &
		"101011100000110101" &
		"00000000000000000000" &
		"011001011011110" &
		"00000000000000000000" &
		"011011110001110111" &
		"00000000000000000000" &
		"1011101101011010" &
		"00000000000000000000" &
		"101110000111101111" &
		"00000000000000000000" &
		"111110001111000110" &
		"00000000000000000000" &
		"01111101111110001" &
		"00000000000000000000" &
		"001010100011100010" &
		"00000000000000000000" &
		"10111000010001000" &
		"00000000000000000000" &
		"101110111111110111" &
		"00000000000000000000" &
		"1010010010000110" &
		"00000000000000000000" &
		"001011111111110" &
		"00000000000000000000" &
		"10110101010110101" &
		"00000000000000000000" &
		"1011001110011" &
		"00000000000000000000" &
		"1010000100100110" &
		"00000000000000000000" &
		"111000111010001110" &
		"00000000000000000000" &
		"1010100010110110" &
		"00000000000000000000" &
		"011001101110101101" &
		"00000000000000000000" &
		"0110110100101000" &
		"00000000000000000000" &
		"0111010000110101" &
		"00000000000000000000" &
		"101111010001110" &
		"00000000000000000000" &
		"1111101001001111" &
		"00000000000000000000" &
		"00111111111000111" &
		"00000000000000000000" &
		"1110110111110000" &
		"00000000000000000000" &
		"11100010110110110" &
		"00000000000000000000" &
		"01111111111110000" &
		"00000000000000000000" &
		"111001111110000011" &
		"00000000000000000000" &
		"111000110101111" &
		"00000000000000000000" &
		"10101110010010110" &
		"00000000000000000000" &
		"11111110111101101" &
		"00000000000000000000" &
		"001110011001010100" &
		"00000000000000000000" &
		"111110000111100001" &
		"00000000000000000000" &
		"111010101110010011" &
		"00000000000000000000" &
		"11100111010101000" &
		"00000000000000000000" &
		"1110011011111011" &
		"00000000000000000000" &
		"011110100010001110" &
		"00000000000000000000" &
		"101001011111" &
		"00000000000000000000" &
		"011010000011111000" &
		"00000000000000000000" &
		"00110010101110" &
		"00000000000000000000" &
		"10111111011001101" &
		"00000000000000000000" &
		"111100100001110000" &
		"00000000000000000000" &
		"00111110101101110" &
		"00000000000000000000" &
		"0011010000101" &
		"00000000000000000000" &
		"01100000010101" &
		"00000000000000000000" &
		"1111100000101111" &
		"00000000000000000000" &
		"0111110111000011" &
		"00000000000000000000" &
		"001100111111001110" &
		"00000000000000000000" &
		"10100001111111110" &
		"00000000000000000000" &
		"001011110011010010" &
		"00000000000000000000" &
		"10110101110" &
		"00000000000000000000" &
		"1110000111010011" &
		"00000000000000000000" &
		"101000000010110100" &
		"00000000000000000000" &
		"101011001011111100" &
		"00000000000000000000" &
		"111001011101010001" &
		"00000000000000000000" &
		"10101101100101110" &
		"00000000000000000000" &
		"101101000100010" &
		"00000000000000000000" &
		"0010101011101110" &
		"00000000000000000000" &
		"0010101100111000" &
		"00000000000000000000" &
		"001110011110101100" &
		"00000000000000000000" &
		"111110101111110110" &
		"00000000000000000000" &
		"101001111010110001" &
		"00000000000000000000" &
		"101100000011111000" &
		"00000000000000000000" &
		"111111101101100010" &
		"00000000000000000000" &
		"111100010000010111" &
		"00000000000000000000" &
		"01101001101101100" &
		"00000000000000000000" &
		"001101101010010100" &
		"00000000000000000000" &
		"011001110101010101" &
		"00000000000000000000" &
		"011001010100101001" &
		"00000000000000000000" &
		"011011111111110100" &
		"00000000000000000000" &
		"001111101101111000" &
		"00000000000000000000" &
		"01100110010000101" &
		"00000000000000000000" &
		"00111110111110011" &
		"00000000000000000000" &
		"011010111011010100" &
		"00000000000000000000" &
		"001000010101011100" &
		"00000000000000000000" &
		"111100110001011001" &
		"00000000000000000000" &
		"011111111011011" &
		"00000000000000000000" &
		"011010100111011110" &
		"00000000000000000000" &
		"011000011010010" &
		"00000000000000000000" &
		"1010100010001111" &
		"00000000000000000000" &
		"101100000000001110" &
		"00000000000000000000" &
		"101101011101001100" &
		"00000000000000000000" &
		"11101100110001111" &
		"00000000000000000000" &
		"1011110000001111" &
		"00000000000000000000" &
		"1011001001110111" &
		"00000000000000000000" &
		"001000001110101010" &
		"00000000000000000000" &
		"011010000100000" &
		"00000000000000000000" &
		"11110101010" &
		"00000000000000000000" &
		"01101010011110110" &
		"00000000000000000000" &
		"11111000011101000" &
		"00000000000000000000" &
		"0010100011100001" &
		"00000000000000000000" &
		"10100000110100010" &
		"00000000000000000000" &
		"01111110010011001" &
		"00000000000000000000" &
		"101100010001100000" &
		"00000000000000000000" &
		"111000010001000111" &
		"00000000000000000000" &
		"001100000111000100" &
		"00000000000000000000" &
		"111000101011001001" &
		"00000000000000000000" &
		"01111100110011000" &
		"00000000000000000000" &
		"111000110011100011" &
		"00000000000000000000" &
		"011110101110000111" &
		"00000000000000000000" &
		"011110111111101001" &
		"00000000000000000000" &
		"001000111011010111" &
		"00000000000000000000" &
		"101110011001001100" &
		"00000000000000000000" &
		"111100011001001000" &
		"00000000000000000000" &
		"001100000001100" &
		"00000000000000000000" &
		"001001000110010000" &
		"00000000000000000000" &
		"111001101010001010" &
		"00000000000000000000" &
		"1110111000110011" &
		"00000000000000000000" &
		"011100101111100011" &
		"00000000000000000000" &
		"11111000010000001" &
		"00000000000000000000" &
		"10101101011100111" &
		"00000000000000000000" &
		"0111111010000000" &
		"00000000000000000000" &
		"0110001111000101" &
		"00000000000000000000" &
		"101010010110010111" &
		"00000000000000000000" &
		"00100000001110011" &
		"00000000000000000000" &
		"011101001100011111" &
		"00000000000000000000" &
		"00100000110110100" &
		"00000000000000000000" &
		"111010100100011110" &
		"00000000000000000000" &
		"1011010010000000" &
		"00000000000000000000" &
		"111101111011011111" &
		"00000000000000000000" &
		"01101000101001" &
		"00000000000000000000" &
		"11100111000101111" &
		"00000000000000000000" &
		"1010100000100" &
		"00000000000000000000" &
		"111010000010000110" &
		"00000000000000000000" &
		"001011011010110011" &
		"00000000000000000000" &
		"01111101010000010" &
		"00000000000000000000" &
		"111110010111011010" &
		"00000000000000000000" &
		"111001110001101101" &
		"00000000000000000000" &
		"111110100110000010" &
		"00000000000000000000" &
		"101110111000111111" &
		"00000000000000000000" &
		"111001010101000011" &
		"00000000000000000000" &
		"011010111110110100" &
		"00000000000000000000" &
		"011010101110001011" &
		"00000000000000000000" &
		"011000011100100010" &
		"00000000000000000000" &
		"10111010111111101" &
		"00000000000000000000" &
		"00111100001000001" &
		"00000000000000000000" &
		"001011111101101111" &
		"00000000000000000000" &
		"011011001000010101" &
		"00000000000000000000" &
		"0010101000010110" &
		"00000000000000000000" &
		"01100110100101010" &
		"00000000000000000000" &
		"0010110110010101" &
		"00000000000000000000" &
		"0010101110000111" &
		"00000000000000000000" &
		"10110001000101110" &
		"00000000000000000000" &
		"111010001010011011" &
		"00000000000000000000" &
		"001101100011110111" &
		"00000000000000000000" &
		"001001001000010010" &
		"00000000000000000000" &
		"011100101010000" &
		"00000000000000000000" &
		"101000011100100110" &
		"00000000000000000000" &
		"101011101001111000" &
		"00000000000000000000" &
		"00111001110001011" &
		"00000000000000000000" &
		"00111100100000000" &
		"00000000000000000000" &
		"11110011110111101" &
		"00000000000000000000" &
		"111010110010000001" &
		"00000000000000000000" &
		"101111110001101010" &
		"00000000000000000000" &
		"111110010010000001" &
		"00000000000000000000" &
		"011000100001111011" &
		"00000000000000000000" &
		"001111101101111110" &
		"00000000000000000000" &
		"001000110111101010" &
		"00000000000000000000" &
		"01101001111011010" &
		"00000000000000000000" &
		"001000001010000000" &
		"00000000000000000000" &
		"111111101110110110" &
		"00000000000000000000" &
		"001000100000011110" &
		"00000000000000000000" &
		"00100100001011100" &
		"00000000000000000000" &
		"0010010001000111" &
		"00000000000000000000" &
		"01110101010011101" &
		"00000000000000000000" &
		"0011111100001001" &
		"00000000000000000000" &
		"111101100010100001" &
		"00000000000000000000" &
		"101010101111011000" &
		"00000000000000000000" &
		"11110100010110000" &
		"00000000000000000000" &
		"111011101000110000" &
		"00000000000000000000" &
		"01100100011111110" &
		"00000000000000000000" &
		"101110101100110000" &
		"00000000000000000000" &
		"001001100010101001" &
		"00000000000000000000" &
		"011111000001010011" &
		"00000000000000000000" &
		"00111000010100101" &
		"00000000000000000000" ;

    -- Channel 2 -> MEM[1] -> 162
    -- Channel 1 -> MEM[2] -> 75

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (
				42095 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				45496 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				12175 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				56445 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				40193 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				35969 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				15369 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				30078 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				9440 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				52689 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				53731 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				32459 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				54649 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				16070 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				21251 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				12660 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				64789 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				9443 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				55107 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				435 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				45808 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				16138 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				25633 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				42763 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				23029 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				28525 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				62610 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				3136 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				1072 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				19049 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				64360 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				41854 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				21137 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				35949 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				30284 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				1445 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				24273 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				39625 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				5499 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				31106 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				33251 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				44154 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				6919 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				31982 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				54486 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				2464 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				20275 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				33920 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				37045 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				53469 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				36081 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				50448 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				38133 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				6772 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				26888 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				12351 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				62900 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				62856 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				11791 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				763 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				38489 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				8934 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				51084 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				37686 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				8509 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				13165 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				53690 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				35891 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				19911 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				20292 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				28640 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				11537 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				44291 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				46031 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				17981 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				37401 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				30455 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				19962 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				37022 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				18917 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				39632 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				36172 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				29467 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				18889 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				20910 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				18179 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				13419 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				20768 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				56288 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				35162 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				47756 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				62635 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				14994 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				7360 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				57800 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				18994 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				28553 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				5672 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				5121 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				11463 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				4948 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				52621 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				22704 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				11087 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				50481 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				4539 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				10775 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				59794 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				2799 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				52424 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				27510 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				24586 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				4102 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				84 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				23229 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				47180 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				39834 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				30415 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				6698 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				52224 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				11487 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				41938 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				37697 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				43240 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				23841 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				44423 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				50904 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				47971 => STD_LOGIC_VECTOR(to_unsigned(190, 8)),
				46252 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				50666 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				58012 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				18667 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				48224 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				9974 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				2438 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				1579 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				24173 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				33739 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				18177 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				14821 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				24146 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				18692 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				9287 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				4476 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				60388 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				63056 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				46605 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				1463 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				16492 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				54281 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				32416 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				27291 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				41615 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				646 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				21232 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				27055 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				56990 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				16132 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				15820 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				6134 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				26447 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				26557 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				10957 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				41847 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				44084 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				28209 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				20488 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				14796 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				30408 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				46559 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				7776 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				63053 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				43139 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				28343 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				35472 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				15242 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				58239 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				3309 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				20606 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				10838 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				31332 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				22002 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				20816 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				25093 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				25018 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				59307 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				13162 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				43986 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				11459 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				62089 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				53414 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				15587 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				23043 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				24310 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				15035 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				28684 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				59058 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				34436 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				59363 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				43269 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				59582 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				19683 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				33719 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				17319 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				2972 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				41784 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				16817 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				23575 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				15108 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				19881 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				2822 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				11661 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				21253 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				39246 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				16877 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				30915 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				63986 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				15550 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				10073 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				43989 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				53332 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				29845 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				63832 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				63162 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				8548 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				47090 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				8941 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				9492 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				53697 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				13946 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				16969 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				62665 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				17942 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				22247 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				21398 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				35516 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				45632 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				20888 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				36909 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				34111 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				27233 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30281 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				39307 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				602 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				3023 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				38089 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				10349 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				11777 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				52879 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				9588 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				16572 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				16675 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				32748 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				38165 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				1319 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				876 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				2734 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				7906 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				59480 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				28574 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				36206 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				64219 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				47503 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				9058 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				51939 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				27184 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				64064 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				64343 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				36840 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				4274 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				13305 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				25284 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				56389 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				32375 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				23143 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				28201 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				15480 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				59713 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				46528 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				59898 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				1889 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				21317 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				48264 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				44053 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				3121 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				29025 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				19511 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				62622 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				35702 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				39783 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				47080 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				61258 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				42396 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				1154 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				54315 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				24739 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				24557 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				15326 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				30649 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				61792 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				12474 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				30472 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				25024 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				62347 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				1122 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				52728 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				1945 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				34144 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				26837 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				53703 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				55335 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				164 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				41347 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				49330 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				277 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				6738 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				36521 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				25266 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				4983 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				48244 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				54731 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				30703 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				18990 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				37740 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				41600 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				58932 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20248 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				45324 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				30101 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				14050 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				20705 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				49844 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				36441 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				46314 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				55650 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				64641 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				34818 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				511 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				32118 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				51002 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				19780 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				13770 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				15506 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				63071 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				688 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				23137 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				55006 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				16256 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				43451 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				45400 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				4205 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				53263 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				62871 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				1071 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				63347 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				41994 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				5946 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				2668 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41796 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				55790 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				62895 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				46327 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				24936 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				48921 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				5881 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				38817 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				53917 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				7650 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				9674 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				5056 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				23336 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				52687 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				54277 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				16208 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				6166 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				24225 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				54381 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				24122 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				48058 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				10369 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				37785 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				59748 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				11660 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				17599 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				12273 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				39042 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				28049 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				20278 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				36708 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				43605 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				14317 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				4843 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				40040 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				61215 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				62630 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				54613 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				21932 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				51409 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				36116 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				23636 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				3256 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				32204 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				64321 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				25984 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				29842 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				58407 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				63659 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				1844 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				48573 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				17503 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				21449 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				42605 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				43551 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				63815 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				43116 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				58279 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				37281 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				54173 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				41787 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				30755 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				62754 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				55305 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				10260 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				43980 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				35417 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				229 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				50437 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				27886 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				6049 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				39157 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				16256 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				4375 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				31505 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				29081 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				13400 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				16080 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				55205 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				55309 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				6168 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				53140 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				34579 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				19411 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				33969 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				21430 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				22888 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				38165 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				49003 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				34561 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				38832 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				6196 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				7135 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				12738 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				1112 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				27945 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				28270 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				22123 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				1626 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				46457 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				47985 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				54967 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				7734 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				62062 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				8315 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				45028 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				49422 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				58770 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				52084 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				42216 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				3601 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				23724 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				39671 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				51057 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				13936 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				58091 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				29559 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				14571 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				21735 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				58210 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				29857 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				11938 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				28003 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				14883 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				41840 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				10017 => STD_LOGIC_VECTOR(to_unsigned(200, 8)),
				42114 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				11374 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				35838 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				21991 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				2246 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				42592 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				26268 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				46305 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				18803 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				14797 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				55039 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				25229 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				2138 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				14253 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				45933 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				18774 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				57424 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				49754 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				51460 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				34082 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				8491 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				62216 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				53280 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				18438 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				50433 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				48536 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				51624 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				61402 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				41873 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				34034 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				40506 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				9562 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				10900 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				53098 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				5914 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				63014 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				59768 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				23136 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				43003 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				26765 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				48938 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				27328 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				14970 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				828 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				12322 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				13514 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				45029 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				25371 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				6348 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				6205 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				41860 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				16352 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				20861 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				64686 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				43688 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				59781 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				43829 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				22572 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				27383 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				63813 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				48675 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				11395 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				34802 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				5395 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				43921 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				7956 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				39852 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				61604 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				42065 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				43181 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				23129 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				16516 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				1771 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				64854 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				39248 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				1017 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				38211 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				27133 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				29747 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				1963 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				56643 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				30833 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				55317 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				8828 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				54860 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				14624 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				29722 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				15596 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				442 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				40587 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				36151 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				62241 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				28926 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				46034 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				6710 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				33762 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				30862 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				60184 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				37543 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				36591 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				13756 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				14789 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				12854 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				28910 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				6092 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				52513 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				62776 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				37727 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				64706 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				49848 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				37242 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				14658 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				60337 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				57094 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				38999 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				34621 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				21879 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				47704 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				28473 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				54504 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				50581 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				47918 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				33050 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				29067 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				967 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				41554 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				38271 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				62852 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				20022 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				62041 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				38989 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				34080 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				10133 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				45364 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				55314 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				54578 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				3762 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				8399 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				13192 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				1733 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				13634 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				40453 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				36258 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				9861 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				33471 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				59991 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				24255 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				55409 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				52519 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				13681 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				9179 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				32981 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				37890 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				11280 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				31469 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				24984 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				24231 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				11772 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				54395 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				18718 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				18383 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				41299 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				33451 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				48958 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				5469 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				44020 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				23085 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				16606 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				58216 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				56768 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				20981 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				41114 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				53591 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				9022 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				6924 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				45358 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				18069 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				58362 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				10281 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				24562 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				25884 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				17406 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				52881 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				57321 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				11093 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				52569 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				50739 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				37836 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				10202 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				51676 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				48806 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				26764 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				42605 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				57374 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				40121 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				39662 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				48206 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				55890 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				36710 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				54273 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				32942 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				35015 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				40964 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				43194 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				21568 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				61264 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				8666 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				13337 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				23378 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				2343 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				39742 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				42120 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				8633 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				41886 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				43658 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				5664 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				21043 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				3309 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				34364 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				51447 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				10382 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				2778 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				44386 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				23244 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				37791 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				54114 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				47743 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				3307 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				57625 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				18028 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				52923 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				62650 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				9450 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				26508 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				41012 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				46439 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				62640 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				52184 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				24037 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				42760 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				60471 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				63604 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				52012 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				18896 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				5741 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				10556 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				35955 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				5854 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				48416 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				34273 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				42484 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				31832 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				38895 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				60279 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				51570 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				2537 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				47862 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				19449 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				6560 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				43128 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				284 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				5392 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				53067 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				33842 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				60342 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				18648 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				35463 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				20779 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				62651 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				51948 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				19129 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				61103 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				30279 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				50829 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				55357 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				46710 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				36280 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				1763 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				18332 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				23465 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				17746 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				58689 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				35000 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				23342 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				40659 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				8546 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				34492 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				26553 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				49590 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				48783 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				62087 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				7282 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				64214 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				265 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				58704 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				17121 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				15768 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				32576 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				20111 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				28882 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				19694 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				49598 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				9998 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				34663 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				3986 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				23917 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				62120 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				28443 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				62690 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				39916 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				37870 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				30594 => STD_LOGIC_VECTOR(to_unsigned(223, 8)),
				42136 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				11929 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				45856 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				36856 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				20645 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				27312 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				24628 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				42107 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				35612 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				51685 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				19008 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				48929 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				7728 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				42852 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				21436 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				42234 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				3415 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				20992 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				18220 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				57437 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				58784 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				47400 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				15599 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				58450 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				8040 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				9443 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				61628 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				20291 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				46227 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				13366 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				47157 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				4830 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				48247 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				15194 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				57839 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				58310 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				31729 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				43234 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				28808 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				61431 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				9350 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				6142 => STD_LOGIC_VECTOR(to_unsigned(162, 8)),
				27317 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				1651 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				8486 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				36494 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				10422 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				39853 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				11560 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				13365 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				7822 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				14927 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				32711 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				11760 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				17846 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				32752 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				40835 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				4527 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				23702 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				32237 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				58964 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				57825 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				43923 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				20136 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				9979 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				59534 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				607 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				41208 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				3246 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				32461 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				51312 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				32110 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				1669 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				2069 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				14383 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				15811 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				53198 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				17406 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				48338 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				430 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				8659 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				32948 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				45820 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				38737 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				23342 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				6690 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				10990 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				11064 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				59308 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				60406 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				40625 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				49400 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				64354 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				50199 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				21356 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				55956 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				40277 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				38185 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				49140 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				64376 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				19589 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				32243 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				44756 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				34140 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				52313 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				8155 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				43486 => STD_LOGIC_VECTOR(to_unsigned(77, 8)),
				4306 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				10383 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				49166 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				55116 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				22927 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				15375 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				12919 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				33706 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				5152 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				426 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				21750 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				28904 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				10465 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				16802 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				31897 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				50272 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				33863 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				49604 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				35529 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				31128 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				36067 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				60295 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				61417 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				36567 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				58956 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				50760 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				6156 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				37264 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				39562 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				11827 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				52195 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				28801 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				23271 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				16000 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				9157 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				42391 => STD_LOGIC_VECTOR(to_unsigned(5, 8)),
				16499 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				54047 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				16820 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				43294 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				13440 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				57055 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				2601 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				20015 => STD_LOGIC_VECTOR(to_unsigned(43, 8)),
				1284 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				41094 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				46771 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				31362 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				58842 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				40045 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				59778 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				60991 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				38211 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				44980 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				43915 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				34594 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				30205 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				30785 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				49007 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				45589 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				10774 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				19754 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				11669 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				11143 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				25134 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				41627 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				55543 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				37394 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				6480 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				34598 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				47736 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				29579 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				30976 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				26557 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				44161 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				64618 => STD_LOGIC_VECTOR(to_unsigned(50, 8)),
				58497 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				34939 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				64382 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				36330 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				21466 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				33408 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				64438 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				34846 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				18524 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				9287 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				27293 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				16137 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				55457 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				43992 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				26800 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				47664 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				18686 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				60208 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				39081 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				61523 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				28837 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),

                              
                                
                                OTHERS => "00000000"-- (OTHERS => '0')
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
            END IF;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        -- wait for 10000 ns;
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        WAIT UNTIL tb_start = '1';
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  62
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  235
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  235
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  132
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  235
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  70
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  235
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  139
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  235
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  139
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  139
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  126
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  116
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  116
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  34
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  49
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  127
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  245
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  219
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  55
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  88
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  222
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  71
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  106
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  58
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  232
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  209
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  209
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  209
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  209
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  46
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  46
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  66
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  66
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  66
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  117
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  66
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  66
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  190
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  192
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  5
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  122
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  235
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  98
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  194
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  51
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  51
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  51
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  3
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(242, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  242
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  251
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  251
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  185
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  185
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(190, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  190
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  206
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  206
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  206
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  206
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  83
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  148
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  148
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  56
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  17
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  56
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  56
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  161
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  161
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  161
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  214
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  241
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  241
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  173
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  173
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  32
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  116
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  106
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  206
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  18
        ASSERT tb_z1 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  206
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  206
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  77
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  159
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  93
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  84
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  93
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  192
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  172
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  11
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  11
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  11
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  203
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  203
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  45
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  45
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  45
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  180
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  186
        ASSERT tb_z3 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  180
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  180
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  165
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  165
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  165
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  26
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  241
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  191
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  152
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  222
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  38
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  222
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  38
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  226
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  195
        ASSERT tb_z3 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  226
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  226
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  77
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  206
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  206
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  60
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  178
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  60
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  178
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  67
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  2
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  2
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  234
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  202
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  198
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  202
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  198
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  254
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  254
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  41
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  168
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  168
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  191
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  33
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  126
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  126
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  24
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  90
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  24
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  130
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  130
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  50
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  50
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  37
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  98
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  98
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  112
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  28
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  112
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  28
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  131
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  47
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  47
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  61
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  47
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  192
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  38
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  153
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  123
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  144
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  43
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  43
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  43
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  43
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  43
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  54
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  54
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  169
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  63
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  63
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  43
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  16
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  16
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  194
        ASSERT tb_z3 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  16
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  191
        ASSERT tb_z3 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  16
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  191
        ASSERT tb_z3 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  141
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  191
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  47
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  136
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  136
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  136
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  195
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  136
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  44
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  136
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  85
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  155
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  240
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  188
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  188
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  47
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  188
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  47
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  57
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  57
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  5
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  57
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  5
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  57
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  57
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  118
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  118
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  118
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  137
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  23
        ASSERT tb_z1 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  137
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  92
        ASSERT tb_z1 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  137
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  137
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  229
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  177
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  229
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  212
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  87
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  31
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  67
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  67
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  5
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  5
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  5
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  152
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  57
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  67
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  67
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  67
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  67
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  67
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  215
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  142
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  94
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  250
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  250
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  166
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  71
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  71
        ASSERT tb_z1 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  189
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  71
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  136
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  86
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  86
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  251
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  211
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  211
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  212
        ASSERT tb_z3 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  96
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  96
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  96
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  154
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  96
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  154
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  5
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  82
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  5
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  5
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  171
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  77
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  148
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  148
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(200, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  200
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(200, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  200
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(200, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  200
        ASSERT tb_z1 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  144
        ASSERT tb_z2 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  53
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(200, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  200
        ASSERT tb_z1 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  144
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(200, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  200
        ASSERT tb_z1 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  144
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  144
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  155
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  23
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  88
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  88
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  88
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  185
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  85
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  88
        ASSERT tb_z3 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  85
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  85
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(150, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  150
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  65
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  99
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  99
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  205
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  99
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  143
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  2
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  2
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  2
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  253
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  164
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  42
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  42
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  116
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  167
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  116
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  167
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  34
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  34
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  56
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  149
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  209
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  60
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  95
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  30
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  30
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  196
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  30
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  34
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  30
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  30
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  131
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  131
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  110
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  84
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  55
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  55
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  156
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  80
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  30
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  30
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  89
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  30
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  165
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  30
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  30
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  182
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  11
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  11
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  153
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  153
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  50
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  145
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  50
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  145
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  145
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  204
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  89
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  89
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  89
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  162
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  162
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  167
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  236
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  104
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  59
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  53
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  74
        ASSERT tb_z3 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  53
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  53
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  131
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  130
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  130
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  193
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  244
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  244
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  244
        ASSERT tb_z3 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  156
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  74
        ASSERT tb_z3 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  156
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  74
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  74
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  175
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  36
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  120
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  3
        ASSERT tb_z2 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  232
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  3
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  3
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  229
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  229
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  92
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  229
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  100
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  100
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  174
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  19
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  76
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  76
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  234
        ASSERT tb_z1 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  76
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  159
        ASSERT tb_z1 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  76
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  159
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  77
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  77
        ASSERT tb_z1 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  156
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  253
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  77
        ASSERT tb_z1 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  156
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  77
        ASSERT tb_z1 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  156
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  77
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  128
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  114
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  39
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  141
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  141
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  141
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  74
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  74
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  163
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  163
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  94
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  94
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  94
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  93
        ASSERT tb_z1 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  50
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  93
        ASSERT tb_z1 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  2
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  93
        ASSERT tb_z1 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  64
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  64
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  122
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  64
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  64
        ASSERT tb_z2 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  218
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  64
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  121
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  162
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  231
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  174
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  174
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  174
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  153
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  174
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  153
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  153
        ASSERT tb_z1 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  20
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  20
        ASSERT tb_z2 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  172
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  20
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  223
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  166
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  166
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  192
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  162
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  162
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  83
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  83
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  9
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  9
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  9
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  69
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  162
        ASSERT tb_z3 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  69
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  69
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  191
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  119
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  32
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  104
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  149
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  156
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  156
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  162
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  162
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  223
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  247
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  170
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  170
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  170
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  170
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  117
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  117
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  220
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  192
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  170
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  164
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(223, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  223
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  231
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  203
        ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  231
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  203
        ASSERT tb_z3 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  231
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  203
        ASSERT tb_z3 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  197
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  197
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  197
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  197
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  197
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  85
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  85
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  41
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  91
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  127
        ASSERT tb_z2 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  91
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  91
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  44
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  99
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  53
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  53
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  53
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(134, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  134
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  53
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  45
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  45
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  116
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  173
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  79
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(162, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  162
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  72
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  130
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  107
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  54
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  246
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  62
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  19
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  33
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  33
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  33
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  4
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  253
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  210
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  147
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  23
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  117
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  215
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  48
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  26
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  21
        ASSERT tb_z1 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  26
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  21
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  155
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(77, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  77
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  219
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  219
        ASSERT tb_z3 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  52
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  122
        ASSERT tb_z3 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  52
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  249
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  52
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  52
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  52
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  115
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  115
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  115
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  115
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  85
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  85
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  231
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  47
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  237
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  47
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  47
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  31
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  220
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  191
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  220
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  191
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  191
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  89
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  59
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  59
        ASSERT tb_z2 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  5
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  59
        ASSERT tb_z2 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  5
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  5
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  5
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(5, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  5
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  212
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  17
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  17
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(43, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  43
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  119
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  119
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  4
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  225
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  102
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  252
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  14
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  106
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  214
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  198
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  95
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  161
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  93
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  119
        ASSERT tb_z1 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  65
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  252
        ASSERT tb_z1 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  65
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  65
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  174
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  174
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  49
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  115
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  66
        ASSERT tb_z1 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  36
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  66
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(50, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  50
        ASSERT tb_z3 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  53
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  121
        ASSERT tb_z3 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  53
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  121
        ASSERT tb_z3 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  69
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  112
        ASSERT tb_z2 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  121
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  121
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  218
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  218
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  218
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  218
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        
        ASSERT false REPORT "Simulation Ended! TEST PASSATO ()" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;
