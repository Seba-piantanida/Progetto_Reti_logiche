
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 35015; -- 5 + 3 + 20 + 7   (RST) + (CH2-MEM[1]) + 20 CYCLES + (CH1-MEM[6])
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00110" & 
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000" &
		"00000000000000000000" &
		"0000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"00000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000" &
		"00000000000000000000" &
		"00000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" &
		"0000000000000000" &
		"00000000000000000000" &
		"000000000000000000" &
		"00000000000000000000" ;

    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000" & 
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111" &
		"00000000000000000000" &
		"1111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"11111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111" &
		"00000000000000000000" &
		"11111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" &
		"1111111111111111" &
		"00000000000000000000" &
		"111111111111111111" &
		"00000000000000000000" ;

    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000" & 
		"0010110001001111" &
		"00000000000000000000" &
		"101111010101001000" &
		"00000000000000000000" &
		"001011110110" &
		"00000000000000000000" &
		"00101100010101000" &
		"00000000000000000000" &
		"011100000010010000" &
		"00000000000000000000" &
		"0110100111000010" &
		"00000000000000000000" &
		"001100010001010011" &
		"00000000000000000000" &
		"101001111110000111" &
		"00000000000000000000" &
		"10111000010000101" &
		"00000000000000000000" &
		"101011011111010001" &
		"00000000000000000000" &
		"001110000110001000" &
		"00000000000000000000" &
		"00111110010101011" &
		"00000000000000000000" &
		"111001000000011100" &
		"00000000000000000000" &
		"101000001100000001" &
		"00000000000000000000" &
		"11101011101110" &
		"00000000000000000000" &
		"01111100011111001" &
		"00000000000000000000" &
		"11111011100010000" &
		"00000000000000000000" &
		"1011101101011100" &
		"00000000000000000000" &
		"11100000001110111" &
		"00000000000000000000" &
		"011010011011100111" &
		"00000000000000000000" &
		"11110000000101100" &
		"00000000000000000000" &
		"10110111010100" &
		"00000000000000000000" &
		"111101010111011" &
		"00000000000000000000" &
		"0011011110000110" &
		"00000000000000000000" &
		"11111111010101110" &
		"00000000000000000000" &
		"0110011001011" &
		"00000000000000000000" &
		"011010011001011000" &
		"00000000000000000000" &
		"00101011100001001" &
		"00000000000000000000" &
		"111001100111001011" &
		"00000000000000000000" &
		"111110011111101100" &
		"00000000000000000000" &
		"101001011000101011" &
		"00000000000000000000" &
		"00100000001001111" &
		"00000000000000000000" &
		"01100011010110011" &
		"00000000000000000000" &
		"111001100010110" &
		"00000000000000000000" &
		"1011001000000011" &
		"00000000000000000000" &
		"111101000111100100" &
		"00000000000000000000" &
		"0111010011110111" &
		"00000000000000000000" &
		"11110010010100000" &
		"00000000000000000000" &
		"11101000110000111" &
		"00000000000000000000" &
		"00100000101111010" &
		"00000000000000000000" &
		"011010110010000" &
		"00000000000000000000" &
		"11101101011110" &
		"00000000000000000000" &
		"011000111000001010" &
		"00000000000000000000" &
		"011100010010101010" &
		"00000000000000000000" &
		"0110100001111" &
		"00000000000000000000" &
		"011000111101101001" &
		"00000000000000000000" &
		"00110010010101011" &
		"00000000000000000000" &
		"101011001" &
		"00000000000000000000" &
		"01101010011111100" &
		"00000000000000000000" &
		"01111111101011110" &
		"00000000000000000000" &
		"101100101110010001" &
		"00000000000000000000" &
		"101110011110001110" &
		"00000000000000000000" &
		"11111100100001111" &
		"00000000000000000000" &
		"1111010000100100" &
		"00000000000000000000" &
		"111001001111110111" &
		"00000000000000000000" &
		"10100110011001" &
		"00000000000000000000" &
		"00111010011000001" &
		"00000000000000000000" &
		"001100010010000011" &
		"00000000000000000000" &
		"111101101110011101" &
		"00000000000000000000" &
		"001010101110010" &
		"00000000000000000000" &
		"00110100011110110" &
		"00000000000000000000" &
		"011100010011111011" &
		"00000000000000000000" &
		"111001001110111001" &
		"00000000000000000000" &
		"011011111001110001" &
		"00000000000000000000" &
		"1111110011011001" &
		"00000000000000000000" &
		"0110011000101100" &
		"00000000000000000000" &
		"10101110000001010" &
		"00000000000000000000" &
		"00110100110101001" &
		"00000000000000000000" &
		"10110001011100000" &
		"00000000000000000000" &
		"001110111001111" &
		"00000000000000000000" &
		"1111110111101000" &
		"00000000000000000000" &
		"001001101110010001" &
		"00000000000000000000" &
		"10101100111010" &
		"00000000000000000000" &
		"11110101000011100" &
		"00000000000000000000" &
		"1011010101010000" &
		"00000000000000000000" &
		"101000010011010011" &
		"00000000000000000000" &
		"11110011010111011" &
		"00000000000000000000" &
		"0110110010011011" &
		"00000000000000000000" &
		"111110100001101111" &
		"00000000000000000000" &
		"101011111110101100" &
		"00000000000000000000" &
		"011110101001001110" &
		"00000000000000000000" &
		"101100010101111001" &
		"00000000000000000000" &
		"11110111000011110" &
		"00000000000000000000" &
		"01111010011011000" &
		"00000000000000000000" &
		"111011111011000011" &
		"00000000000000000000" &
		"00101000101100101" &
		"00000000000000000000" &
		"101101111110110" &
		"00000000000000000000" &
		"111101110011001000" &
		"00000000000000000000" &
		"101111010110111000" &
		"00000000000000000000" &
		"1111011011011000" &
		"00000000000000000000" &
		"001000101111011000" &
		"00000000000000000000" &
		"001100100100110111" &
		"00000000000000000000" &
		"111100010101001001" &
		"00000000000000000000" &
		"0110011110100010" &
		"00000000000000000000" &
		"011000010010001001" &
		"00000000000000000000" &
		"00101011001101000" &
		"00000000000000000000" &
		"111111011001101001" &
		"00000000000000000000" &
		"10100100001101100" &
		"00000000000000000000" &
		"01111001010001000" &
		"00000000000000000000" &
		"10100000111010111" &
		"00000000000000000000" &
		"10100101001110111" &
		"00000000000000000000" &
		"001110100001000110" &
		"00000000000000000000" &
		"111110001110111" &
		"00000000000000000000" &
		"01111011010100110" &
		"00000000000000000000" &
		"001000100111110111" &
		"00000000000000000000" &
		"10110001011111001" &
		"00000000000000000000" &
		"101110100101010011" &
		"00000000000000000000" &
		"01100001111000111" &
		"00000000000000000000" &
		"011101100100001111" &
		"00000000000000000000" &
		"11101001001101101" &
		"00000000000000000000" &
		"101011101001001011" &
		"00000000000000000000" &
		"00111000011011111" &
		"00000000000000000000" &
		"011000010000010101" &
		"00000000000000000000" &
		"11110000001111" &
		"00000000000000000000" &
		"101001011110010011" &
		"00000000000000000000" &
		"011111110110110011" &
		"00000000000000000000" &
		"11100011100000101" &
		"00000000000000000000" &
		"00101100011111110" &
		"00000000000000000000" &
		"1010111000100" &
		"00000000000000000000" &
		"1010110001111111" &
		"00000000000000000000" &
		"1111011011011" &
		"00000000000000000000" &
		"101100011010000000" &
		"00000000000000000000" &
		"111101100011011100" &
		"00000000000000000000" &
		"00101010000101" &
		"00000000000000000000" &
		"10111110110100101" &
		"00000000000000000000" &
		"01101001111101000" &
		"00000000000000000000" &
		"0011001111001000" &
		"00000000000000000000" &
		"011000001010101000" &
		"00000000000000000000" &
		"001111011110100000" &
		"00000000000000000000" &
		"111110111110101110" &
		"00000000000000000000" &
		"001111110010010101" &
		"00000000000000000000" &
		"011100001010100001" &
		"00000000000000000000" &
		"1111100001101001" &
		"00000000000000000000" &
		"0011100001010011" &
		"00000000000000000000" &
		"111000011110110011" &
		"00000000000000000000" &
		"001100010100010110" &
		"00000000000000000000" &
		"1111010011010010" &
		"00000000000000000000" &
		"011001011010101110" &
		"00000000000000000000" &
		"101100011001" &
		"00000000000000000000" &
		"10101000111111100" &
		"00000000000000000000" &
		"11101101111101110" &
		"00000000000000000000" &
		"011010010110010011" &
		"00000000000000000000" &
		"111100010011101100" &
		"00000000000000000000" &
		"001101010110010111" &
		"00000000000000000000" &
		"001110001101101111" &
		"00000000000000000000" &
		"011010101111100101" &
		"00000000000000000000" &
		"111011100001110101" &
		"00000000000000000000" &
		"111001011000111000" &
		"00000000000000000000" &
		"011111100100110101" &
		"00000000000000000000" &
		"011000101000001110" &
		"00000000000000000000" &
		"00100110000011001" &
		"00000000000000000000" &
		"0011111100011010" &
		"00000000000000000000" &
		"101000001010101101" &
		"00000000000000000000" &
		"101010110010111110" &
		"00000000000000000000" &
		"001100011111011111" &
		"00000000000000000000" &
		"11100101101000111" &
		"00000000000000000000" &
		"011000001001100100" &
		"00000000000000000000" &
		"1111000100111110" &
		"00000000000000000000" &
		"11110000010010111" &
		"00000000000000000000" &
		"11111011101110010" &
		"00000000000000000000" &
		"111101000011111011" &
		"00000000000000000000" &
		"101110001101000111" &
		"00000000000000000000" &
		"011010111110001101" &
		"00000000000000000000" &
		"10111001101110000" &
		"00000000000000000000" &
		"011000101110010110" &
		"00000000000000000000" &
		"011011101101100111" &
		"00000000000000000000" &
		"00100000100001100" &
		"00000000000000000000" &
		"011010100101001110" &
		"00000000000000000000" &
		"101100010000100000" &
		"00000000000000000000" &
		"011101110011000010" &
		"00000000000000000000" &
		"1110001101001100" &
		"00000000000000000000" &
		"111101010010011111" &
		"00000000000000000000" &
		"00110001111110101" &
		"00000000000000000000" &
		"011000111010000101" &
		"00000000000000000000" &
		"111101101001101001" &
		"00000000000000000000" &
		"011110011011100010" &
		"00000000000000000000" &
		"011001010010111001" &
		"00000000000000000000" &
		"111010000111100100" &
		"00000000000000000000" &
		"011100110001100001" &
		"00000000000000000000" &
		"011010001110100" &
		"00000000000000000000" &
		"0111110100111111" &
		"00000000000000000000" &
		"111110001111011010" &
		"00000000000000000000" &
		"1011110111011101" &
		"00000000000000000000" &
		"10101001111111101" &
		"00000000000000000000" &
		"11110111110101011" &
		"00000000000000000000" &
		"0011010101001111" &
		"00000000000000000000" &
		"10100100101001110" &
		"00000000000000000000" &
		"111001111100011" &
		"00000000000000000000" &
		"101111010111111010" &
		"00000000000000000000" &
		"001100010101101010" &
		"00000000000000000000" &
		"111100001101110011" &
		"00000000000000000000" &
		"101010010100010111" &
		"00000000000000000000" &
		"01100001010110101" &
		"00000000000000000000" &
		"10111001101010100" &
		"00000000000000000000" &
		"10101111110010110" &
		"00000000000000000000" &
		"001010101111001101" &
		"00000000000000000000" &
		"00111000010010001" &
		"00000000000000000000" &
		"111011011010010010" &
		"00000000000000000000" &
		"001100111111110011" &
		"00000000000000000000" &
		"11101100010001110" &
		"00000000000000000000" &
		"1010111000110100" &
		"00000000000000000000" &
		"111011010010101101" &
		"00000000000000000000" &
		"001101110101110111" &
		"00000000000000000000" &
		"1111011001111100" &
		"00000000000000000000" &
		"0011100000000" &
		"00000000000000000000" &
		"011100001111001011" &
		"00000000000000000000" &
		"01110010110100001" &
		"00000000000000000000" &
		"1011010011" &
		"00000000000000000000" &
		"101000110111010101" &
		"00000000000000000000" &
		"00110110000101111" &
		"00000000000000000000" &
		"111110000011100010" &
		"00000000000000000000" &
		"001110110100100011" &
		"00000000000000000000" &
		"1110000010010001" &
		"00000000000000000000" &
		"1011101110001110" &
		"00000000000000000000" &
		"00110110001101101" &
		"00000000000000000000" &
		"10111011111001101" &
		"00000000000000000000" &
		"111100101010001110" &
		"00000000000000000000" &
		"001000110011010000" &
		"00000000000000000000" &
		"001111001001111001" &
		"00000000000000000000" &
		"001100000110100010" &
		"00000000000000000000" &
		"011001001100011100" &
		"00000000000000000000" &
		"001111100111101010" &
		"00000000000000000000" &
		"101101011100011100" &
		"00000000000000000000" &
		"111001111011100010" &
		"00000000000000000000" &
		"101001000100001011" &
		"00000000000000000000" &
		"101011101101101010" &
		"00000000000000000000" &
		"11100001001110110" &
		"00000000000000000000" &
		"011001011011101000" &
		"00000000000000000000" &
		"011010101000110100" &
		"00000000000000000000" &
		"0111010010" &
		"00000000000000000000" &
		"001101101100011" &
		"00000000000000000000" &
		"111101111101110001" &
		"00000000000000000000" &
		"00111100010111000" &
		"00000000000000000000" &
		"011100110000" &
		"00000000000000000000" &
		"10100111110110010" &
		"00000000000000000000" &
		"10110111111000000" &
		"00000000000000000000" &
		"01110110111001001" &
		"00000000000000000000" &
		"11111011011001100" &
		"00000000000000000000" &
		"001100110001001100" &
		"00000000000000000000" &
		"11100110011000101" &
		"00000000000000000000" &
		"101010110011011010" &
		"00000000000000000000" &
		"111101011000000101" &
		"00000000000000000000" &
		"101111001100100001" &
		"00000000000000000000" &
		"111101101011101100" &
		"00000000000000000000" &
		"111111101010001001" &
		"00000000000000000000" &
		"1111100101101111" &
		"00000000000000000000" &
		"101111011000110001" &
		"00000000000000000000" &
		"01110100001111110" &
		"00000000000000000000" &
		"11100111010111011" &
		"00000000000000000000" &
		"011011100111" &
		"00000000000000000000" &
		"01101011010010" &
		"00000000000000000000" &
		"001001111111110000" &
		"00000000000000000000" &
		"01110100001010011" &
		"00000000000000000000" &
		"1011010001010001" &
		"00000000000000000000" &
		"10100001010100010" &
		"00000000000000000000" &
		"1010111011001110" &
		"00000000000000000000" &
		"0011101011010100" &
		"00000000000000000000" &
		"001101111100001100" &
		"00000000000000000000" &
		"011110100001010010" &
		"00000000000000000000" &
		"101010011100010011" &
		"00000000000000000000" &
		"101000011001011101" &
		"00000000000000000000" &
		"011100100011011110" &
		"00000000000000000000" &
		"001000110011111100" &
		"00000000000000000000" &
		"0111101110100110" &
		"00000000000000000000" &
		"001001011010010101" &
		"00000000000000000000" &
		"011111011000100111" &
		"00000000000000000000" &
		"111110110000000110" &
		"00000000000000000000" &
		"10100110111011001" &
		"00000000000000000000" &
		"01100001111101011" &
		"00000000000000000000" &
		"101010111000001110" &
		"00000000000000000000" &
		"01100100111000100" &
		"00000000000000000000" &
		"111101010110101000" &
		"00000000000000000000" &
		"101101101100010100" &
		"00000000000000000000" &
		"101001110111110111" &
		"00000000000000000000" &
		"101100110110110110" &
		"00000000000000000000" &
		"011001001111001" &
		"00000000000000000000" &
		"0010101110001111" &
		"00000000000000000000" &
		"1111001011001101" &
		"00000000000000000000" &
		"11111101010011000" &
		"00000000000000000000" &
		"001100011011000000" &
		"00000000000000000000" &
		"10100111000000110" &
		"00000000000000000000" &
		"0011111011100000" &
		"00000000000000000000" &
		"111011110100110011" &
		"00000000000000000000" &
		"001110011000111" &
		"00000000000000000000" &
		"01100111110011000" &
		"00000000000000000000" &
		"10101110000111" &
		"00000000000000000000" &
		"101011001010101001" &
		"00000000000000000000" &
		"10101111001111110" &
		"00000000000000000000" &
		"101001011110101000" &
		"00000000000000000000" &
		"001010010110100011" &
		"00000000000000000000" &
		"011011100011010000" &
		"00000000000000000000" &
		"101001111001100001" &
		"00000000000000000000" &
		"111000001000001101" &
		"00000000000000000000" &
		"101010100010100111" &
		"00000000000000000000" &
		"11110110111001100" &
		"00000000000000000000" &
		"001011011011" &
		"00000000000000000000" &
		"011010001100011000" &
		"00000000000000000000" &
		"11100011111101110" &
		"00000000000000000000" &
		"111101010110101" &
		"00000000000000000000" &
		"0111111011001111" &
		"00000000000000000000" &
		"011110000011010010" &
		"00000000000000000000" &
		"101111001110111100" &
		"00000000000000000000" &
		"01110111001001" &
		"00000000000000000000" &
		"1111000101111000" &
		"00000000000000000000" &
		"011000111110100100" &
		"00000000000000000000" &
		"001110101101011111" &
		"00000000000000000000" &
		"11101010100111" &
		"00000000000000000000" &
		"11110100000111111" &
		"00000000000000000000" &
		"101011100110101001" &
		"00000000000000000000" &
		"011101011110100000" &
		"00000000000000000000" &
		"11111100001100101" &
		"00000000000000000000" &
		"011100110110111000" &
		"00000000000000000000" &
		"011100000100111111" &
		"00000000000000000000" &
		"001100101011001010" &
		"00000000000000000000" &
		"001101001110000100" &
		"00000000000000000000" &
		"0110000100110010" &
		"00000000000000000000" &
		"001011101100100110" &
		"00000000000000000000" &
		"101110001111110" &
		"00000000000000000000" &
		"001000100100000101" &
		"00000000000000000000" &
		"1010010010010010" &
		"00000000000000000000" &
		"011000000001100000" &
		"00000000000000000000" &
		"011000111111111010" &
		"00000000000000000000" &
		"111110001000000100" &
		"00000000000000000000" &
		"001000010000010001" &
		"00000000000000000000" &
		"101101100101111101" &
		"00000000000000000000" &
		"111100000001110011" &
		"00000000000000000000" &
		"101110011000111000" &
		"00000000000000000000" &
		"011011110111110" &
		"00000000000000000000" &
		"111100100000110001" &
		"00000000000000000000" &
		"011011111010110011" &
		"00000000000000000000" &
		"011101010100001001" &
		"00000000000000000000" &
		"011100101001010100" &
		"00000000000000000000" &
		"01100011000101111" &
		"00000000000000000000" &
		"101100100000000011" &
		"00000000000000000000" &
		"10101100000000001" &
		"00000000000000000000" &
		"10101010101011000" &
		"00000000000000000000" &
		"1010101010001111" &
		"00000000000000000000" &
		"011001011001101001" &
		"00000000000000000000" &
		"001001000000011" &
		"00000000000000000000" &
		"10111100110000000" &
		"00000000000000000000" &
		"1110001001011010" &
		"00000000000000000000" &
		"10101111100011110" &
		"00000000000000000000" &
		"1111011100011100" &
		"00000000000000000000" &
		"10101100110101111" &
		"00000000000000000000" &
		"10100010101110001" &
		"00000000000000000000" &
		"111110000100001110" &
		"00000000000000000000" &
		"101101011000111010" &
		"00000000000000000000" &
		"101011101001010000" &
		"00000000000000000000" &
		"011101011110100101" &
		"00000000000000000000" &
		"001001001101000101" &
		"00000000000000000000" &
		"11101111110111000" &
		"00000000000000000000" &
		"001010100011010001" &
		"00000000000000000000" &
		"11110100010101000" &
		"00000000000000000000" &
		"001111000101000101" &
		"00000000000000000000" &
		"001101111010000101" &
		"00000000000000000000" &
		"111110000100100100" &
		"00000000000000000000" &
		"00100000111000111" &
		"00000000000000000000" &
		"111011010001101110" &
		"00000000000000000000" &
		"111000000110000011" &
		"00000000000000000000" &
		"011100110001101111" &
		"00000000000000000000" &
		"011010011111001010" &
		"00000000000000000000" &
		"0111010011110011" &
		"00000000000000000000" &
		"101000100110010101" &
		"00000000000000000000" &
		"011100011010110" &
		"00000000000000000000" &
		"011111101111010010" &
		"00000000000000000000" &
		"01111101001101100" &
		"00000000000000000000" &
		"001110010100011010" &
		"00000000000000000000" &
		"1110101011001010" &
		"00000000000000000000" &
		"001110100000000110" &
		"00000000000000000000" &
		"10101100010011011" &
		"00000000000000000000" &
		"001101110011010100" &
		"00000000000000000000" &
		"1110110001011011" &
		"00000000000000000000" &
		"10101111111110011" &
		"00000000000000000000" &
		"101001101010110101" &
		"00000000000000000000" &
		"00100111001111011" &
		"00000000000000000000" &
		"10111011001110001" &
		"00000000000000000000" &
		"111010111001000010" &
		"00000000000000000000" &
		"01111000010010000" &
		"00000000000000000000" &
		"111110110011100100" &
		"00000000000000000000" &
		"101100001111101" &
		"00000000000000000000" &
		"011011110100111110" &
		"00000000000000000000" &
		"011101001111100001" &
		"00000000000000000000" &
		"0110001111100001" &
		"00000000000000000000" &
		"101111000010010011" &
		"00000000000000000000" &
		"101011011101100000" &
		"00000000000000000000" &
		"10101110010010000" &
		"00000000000000000000" &
		"111011011110111110" &
		"00000000000000000000" &
		"101001101110001001" &
		"00000000000000000000" &
		"001101110010" &
		"00000000000000000000" &
		"1010011000101000" &
		"00000000000000000000" &
		"10100011111101000" &
		"00000000000000000000" &
		"101110011000111011" &
		"00000000000000000000" &
		"10110011111100110" &
		"00000000000000000000" &
		"111010011110101" &
		"00000000000000000000" &
		"101001100110000010" &
		"00000000000000000000" &
		"01100000001010001" &
		"00000000000000000000" &
		"101101111100001001" &
		"00000000000000000000" &
		"0110000111100" &
		"00000000000000000000" &
		"111010111000011110" &
		"00000000000000000000" &
		"01101110" &
		"00000000000000000000" &
		"011011011010010010" &
		"00000000000000000000" &
		"11100011000110010" &
		"00000000000000000000" &
		"111001011100011001" &
		"00000000000000000000" &
		"011111100011101000" &
		"00000000000000000000" &
		"011010101010000001" &
		"00000000000000000000" &
		"1011100100000110" &
		"00000000000000000000" &
		"01110101000001010" &
		"00000000000000000000" &
		"10111101100001011" &
		"00000000000000000000" &
		"0010110110101000" &
		"00000000000000000000" &
		"111101010010000" &
		"00000000000000000000" &
		"111111101111111111" &
		"00000000000000000000" &
		"111111000100010110" &
		"00000000000000000000" &
		"001010100010011110" &
		"00000000000000000000" &
		"101000010011100101" &
		"00000000000000000000" &
		"001101001101011010" &
		"00000000000000000000" &
		"101110011000111100" &
		"00000000000000000000" &
		"01110010001010110" &
		"00000000000000000000" &
		"01110000110111100" &
		"00000000000000000000" &
		"001001100111001001" &
		"00000000000000000000" &
		"111111000111111010" &
		"00000000000000000000" &
		"11110110001100100" &
		"00000000000000000000" &
		"011001111100001100" &
		"00000000000000000000" &
		"00110000110000" &
		"00000000000000000000" &
		"101110001111111000" &
		"00000000000000000000" &
		"101100110011001100" &
		"00000000000000000000" &
		"101000100100000110" &
		"00000000000000000000" &
		"11111001011011001" &
		"00000000000000000000" &
		"10110111010111101" &
		"00000000000000000000" &
		"011111110010101110" &
		"00000000000000000000" &
		"11111100111111000" &
		"00000000000000000000" &
		"101100100001000" &
		"00000000000000000000" &
		"1111100101000101" &
		"00000000000000000000" &
		"10100001100001011" &
		"00000000000000000000" &
		"001001011001101" &
		"00000000000000000000" &
		"101111011111001" &
		"00000000000000000000" &
		"101110110010101011" &
		"00000000000000000000" &
		"00101010111110010" &
		"00000000000000000000" &
		"111110101000101110" &
		"00000000000000000000" &
		"10110001110101000" &
		"00000000000000000000" &
		"001110010010001111" &
		"00000000000000000000" &
		"10101000010111110" &
		"00000000000000000000" &
		"00100010010000101" &
		"00000000000000000000" &
		"001001011101101100" &
		"00000000000000000000" &
		"011000001101011011" &
		"00000000000000000000" &
		"011110111011000001" &
		"00000000000000000000" &
		"01111101011000000" &
		"00000000000000000000" &
		"101101101101001101" &
		"00000000000000000000" &
		"111010110001001100" &
		"00000000000000000000" &
		"11111101011101101" &
		"00000000000000000000" &
		"0110010000001010" &
		"00000000000000000000" &
		"00101001001011" &
		"00000000000000000000" &
		"11111101111100011" &
		"00000000000000000000" &
		"111000110001010101" &
		"00000000000000000000" &
		"001111110011100" &
		"00000000000000000000" &
		"111101000100010110" &
		"00000000000000000000" &
		"001000110011110101" &
		"00000000000000000000" &
		"11110101101101110" &
		"00000000000000000000" &
		"11111111011" &
		"00000000000000000000" &
		"001011011010100000" &
		"00000000000000000000" &
		"11100100101111001" &
		"00000000000000000000" &
		"00101000101110000" &
		"00000000000000000000" &
		"00100100111111100" &
		"00000000000000000000" &
		"10110110110000111" &
		"00000000000000000000" &
		"0110101000010111" &
		"00000000000000000000" &
		"001010101111001011" &
		"00000000000000000000" &
		"001001110101100111" &
		"00000000000000000000" &
		"01111100011000" &
		"00000000000000000000" &
		"101001100111011101" &
		"00000000000000000000" &
		"111011110000001111" &
		"00000000000000000000" &
		"011000101100011000" &
		"00000000000000000000" &
		"111100001000001011" &
		"00000000000000000000" &
		"111110101100111110" &
		"00000000000000000000" &
		"001011101101" &
		"00000000000000000000" &
		"111010011100111" &
		"00000000000000000000" &
		"01110110001100" &
		"00000000000000000000" &
		"0110011001111101" &
		"00000000000000000000" &
		"001111101101001111" &
		"00000000000000000000" &
		"11110010111011000" &
		"00000000000000000000" &
		"011100011111101000" &
		"00000000000000000000" &
		"011100011100001010" &
		"00000000000000000000" &
		"001100111101010100" &
		"00000000000000000000" &
		"01101010100110" &
		"00000000000000000000" &
		"111101011110111001" &
		"00000000000000000000" &
		"0011001100110010" &
		"00000000000000000000" &
		"10100110101000000" &
		"00000000000000000000" &
		"111000010001111100" &
		"00000000000000000000" &
		"001110100000101110" &
		"00000000000000000000" &
		"111111000001110011" &
		"00000000000000000000" &
		"101000000100100" &
		"00000000000000000000" &
		"011000011110101" &
		"00000000000000000000" &
		"00101010001010110" &
		"00000000000000000000" &
		"11110001100100001" &
		"00000000000000000000" &
		"001111011111010000" &
		"00000000000000000000" &
		"001100110110100110" &
		"00000000000000000000" &
		"11110110001101111" &
		"00000000000000000000" &
		"001110110000111100" &
		"00000000000000000000" &
		"011010110010101011" &
		"00000000000000000000" &
		"001101110010011110" &
		"00000000000000000000" &
		"011000100110010101" &
		"00000000000000000000" &
		"001001001101010" &
		"00000000000000000000" &
		"011101100000110011" &
		"00000000000000000000" &
		"1110000010111101" &
		"00000000000000000000" &
		"111010111100101000" &
		"00000000000000000000" &
		"101011111000110101" &
		"00000000000000000000" &
		"111010111101011000" &
		"00000000000000000000" &
		"011110101011100011" &
		"00000000000000000000" &
		"111010100010000101" &
		"00000000000000000000" &
		"011011001110010000" &
		"00000000000000000000" &
		"011100111001100010" &
		"00000000000000000000" &
		"011110011001110000" &
		"00000000000000000000" &
		"011110100011111110" &
		"00000000000000000000" &
		"11110100101101101" &
		"00000000000000000000" &
		"11111101100100001" &
		"00000000000000000000" &
		"101001000001011001" &
		"00000000000000000000" &
		"0011010010110101" &
		"00000000000000000000" &
		"0111011011110110" &
		"00000000000000000000" &
		"001101001111110110" &
		"00000000000000000000" &
		"111010101010010001" &
		"00000000000000000000" &
		"0010110001101110" &
		"00000000000000000000" &
		"00111000110111011" &
		"00000000000000000000" &
		"101110110100001001" &
		"00000000000000000000" &
		"001011100100101110" &
		"00000000000000000000" &
		"1110000001110001" &
		"00000000000000000000" &
		"00111110010111000" &
		"00000000000000000000" &
		"01101111011111000" &
		"00000000000000000000" &
		"10110000011101000" &
		"00000000000000000000" &
		"0110011101110000" &
		"00000000000000000000" &
		"011011010100010000" &
		"00000000000000000000" &
		"101110010100000011" &
		"00000000000000000000" &
		"00111100000111111" &
		"00000000000000000000" &
		"101010010101000001" &
		"00000000000000000000" &
		"11101000010011010" &
		"00000000000000000000" &
		"00111011000101" &
		"00000000000000000000" &
		"001101100011110110" &
		"00000000000000000000" &
		"011111110100001010" &
		"00000000000000000000" &
		"111100011111110100" &
		"00000000000000000000" &
		"011001101100101011" &
		"00000000000000000000" &
		"101011110010110000" &
		"00000000000000000000" &
		"011011010000000011" &
		"00000000000000000000" &
		"01111110011101100" &
		"00000000000000000000" &
		"001110110111100110" &
		"00000000000000000000" &
		"101010100011001" &
		"00000000000000000000" &
		"1011000100000101" &
		"00000000000000000000" &
		"001111100001111010" &
		"00000000000000000000" &
		"1011001001100110" &
		"00000000000000000000" &
		"101111100110001111" &
		"00000000000000000000" &
		"001010001111101000" &
		"00000000000000000000" &
		"01111101111101101" &
		"00000000000000000000" &
		"1011101001100010" &
		"00000000000000000000" &
		"111110100011101101" &
		"00000000000000000000" &
		"011001111110010101" &
		"00000000000000000000" &
		"011001111110111110" &
		"00000000000000000000" &
		"0011010111101011" &
		"00000000000000000000" &
		"101010110000011100" &
		"00000000000000000000" &
		"111010110000011011" &
		"00000000000000000000" &
		"1111000110101010" &
		"00000000000000000000" &
		"0011000100101001" &
		"00000000000000000000" &
		"001000110111010101" &
		"00000000000000000000" &
		"101111110000010111" &
		"00000000000000000000" &
		"011000000110101111" &
		"00000000000000000000" &
		"00111110000100" &
		"00000000000000000000" &
		"101001111110001111" &
		"00000000000000000000" &
		"11111101011011110" &
		"00000000000000000000" &
		"0110100011110011" &
		"00000000000000000000" &
		"00101010100001100" &
		"00000000000000000000" &
		"101111100000000000" &
		"00000000000000000000" &
		"11111100001100" &
		"00000000000000000000" &
		"101111101011111011" &
		"00000000000000000000" &
		"1110101000011110" &
		"00000000000000000000" &
		"00111011101011000" &
		"00000000000000000000" &
		"001010101001101001" &
		"00000000000000000000" &
		"00110011111010101" &
		"00000000000000000000" &
		"101001011011000111" &
		"00000000000000000000" &
		"10110010011001110" &
		"00000000000000000000" &
		"001001110001111100" &
		"00000000000000000000" &
		"1010000111100110" &
		"00000000000000000000" &
		"1111001110100101" &
		"00000000000000000000" &
		"10111101010011001" &
		"00000000000000000000" &
		"101011100010000" &
		"00000000000000000000" &
		"1010100000110101" &
		"00000000000000000000" &
		"001110010001010001" &
		"00000000000000000000" &
		"00101011110011111" &
		"00000000000000000000" &
		"11101000101110001" &
		"00000000000000000000" &
		"101110000101100100" &
		"00000000000000000000" &
		"001110011100111111" &
		"00000000000000000000" &
		"101011011000101001" &
		"00000000000000000000" &
		"011010010111110011" &
		"00000000000000000000" &
		"001100101111110110" &
		"00000000000000000000" &
		"1110111000100011" &
		"00000000000000000000" &
		"1110111111010111" &
		"00000000000000000000" &
		"101011000101" &
		"00000000000000000000" &
		"001111000110010111" &
		"00000000000000000000" &
		"011100010100110011" &
		"00000000000000000000" &
		"11111000010010101" &
		"00000000000000000000" &
		"011111101110101101" &
		"00000000000000000000" &
		"10110100110101101" &
		"00000000000000000000" &
		"011100100010101011" &
		"00000000000000000000" &
		"101001001111111010" &
		"00000000000000000000" &
		"101001111000010" &
		"00000000000000000000" &
		"011000011100001110" &
		"00000000000000000000" &
		"01101000011010101" &
		"00000000000000000000" &
		"001011111001111" &
		"00000000000000000000" &
		"111100110111101100" &
		"00000000000000000000" &
		"011001011111100111" &
		"00000000000000000000" &
		"111111000111101010" &
		"00000000000000000000" &
		"011010110011011111" &
		"00000000000000000000" &
		"111100101010010001" &
		"00000000000000000000" &
		"00111000001001010" &
		"00000000000000000000" &
		"00100111001111" &
		"00000000000000000000" &
		"0111101111011101" &
		"00000000000000000000" &
		"111101101000110011" &
		"00000000000000000000" &
		"01101011011001100" &
		"00000000000000000000" &
		"011101001001011100" &
		"00000000000000000000" &
		"001101100111101100" &
		"00000000000000000000" &
		"011010101001010011" &
		"00000000000000000000" &
		"111000010100000010" &
		"00000000000000000000" &
		"101111000011000" &
		"00000000000000000000" &
		"11110101010100001" &
		"00000000000000000000" &
		"001010001100" &
		"00000000000000000000" &
		"011001100110011100" &
		"00000000000000000000" &
		"111110110110001111" &
		"00000000000000000000" &
		"001010100101111010" &
		"00000000000000000000" &
		"001101011101010000" &
		"00000000000000000000" &
		"101101111110101001" &
		"00000000000000000000" &
		"001101100100101011" &
		"00000000000000000000" &
		"001111011010100111" &
		"00000000000000000000" &
		"11101011110110100" &
		"00000000000000000000" &
		"001011101000000001" &
		"00000000000000000000" &
		"001111000100001010" &
		"00000000000000000000" &
		"0110101010111111" &
		"00000000000000000000" &
		"0010010011010000" &
		"00000000000000000000" &
		"001000100101110" &
		"00000000000000000000" &
		"10110101001010010" &
		"00000000000000000000" &
		"111010001111100101" &
		"00000000000000000000" &
		"111110100110101" &
		"00000000000000000000" &
		"011110001110011010" &
		"00000000000000000000" &
		"10100011001111011" &
		"00000000000000000000" &
		"101000110100001010" &
		"00000000000000000000" &
		"00110010011111000" &
		"00000000000000000000" &
		"101011110101000101" &
		"00000000000000000000" &
		"111000101110010110" &
		"00000000000000000000" &
		"111110101010000" &
		"00000000000000000000" &
		"001100010001111000" &
		"00000000000000000000" &
		"111011010000110100" &
		"00000000000000000000" &
		"001111010000111100" &
		"00000000000000000000" &
		"001010110001000010" &
		"00000000000000000000" &
		"011001010101000011" &
		"00000000000000000000" &
		"011011010001111001" &
		"00000000000000000000" &
		"111111000110101000" &
		"00000000000000000000" &
		"101000110111110000" &
		"00000000000000000000" &
		"0010000101001110" &
		"00000000000000000000" &
		"10110100001100000" &
		"00000000000000000000" &
		"001011110010100101" &
		"00000000000000000000" &
		"0011011110011011" &
		"00000000000000000000" &
		"0111000101001" &
		"00000000000000000000" &
		"111000011011110001" &
		"00000000000000000000" &
		"00100100100111000" &
		"00000000000000000000" &
		"011011010010100011" &
		"00000000000000000000" &
		"011110100000001111" &
		"00000000000000000000" &
		"0011011110111101" &
		"00000000000000000000" &
		"01101010011001111" &
		"00000000000000000000" &
		"01110111001111010" &
		"00000000000000000000" &
		"11100001100011100" &
		"00000000000000000000" &
		"0110110000100000" &
		"00000000000000000000" &
		"011111101000101110" &
		"00000000000000000000" &
		"10110101100110000" &
		"00000000000000000000" &
		"0110100100111001" &
		"00000000000000000000" &
		"01110011111110111" &
		"00000000000000000000" &
		"001100000110110010" &
		"00000000000000000000" &
		"01110011111101010" &
		"00000000000000000000" &
		"001111100110011111" &
		"00000000000000000000" &
		"10111010111001010" &
		"00000000000000000000" &
		"001100010001011111" &
		"00000000000000000000" &
		"111011100010110100" &
		"00000000000000000000" &
		"011011110110101" &
		"00000000000000000000" &
		"01110111101110011" &
		"00000000000000000000" &
		"101001110010011101" &
		"00000000000000000000" &
		"10100111001100001" &
		"00000000000000000000" &
		"011001101010000111" &
		"00000000000000000000" &
		"101100111110001" &
		"00000000000000000000" &
		"11100100000011011" &
		"00000000000000000000" &
		"0110001010010111" &
		"00000000000000000000" &
		"11110111010111011" &
		"00000000000000000000" &
		"01100111110100011" &
		"00000000000000000000" &
		"011010111101001" &
		"00000000000000000000" &
		"001101000000000001" &
		"00000000000000000000" &
		"01101010100110000" &
		"00000000000000000000" &
		"10111111101010101" &
		"00000000000000000000" &
		"101011100000110111" &
		"00000000000000000000" &
		"10111010011111101" &
		"00000000000000000000" &
		"101010111011111011" &
		"00000000000000000000" &
		"10101010110100001" &
		"00000000000000000000" &
		"011111001110000011" &
		"00000000000000000000" &
		"101000000001100001" &
		"00000000000000000000" &
		"011011011010000100" &
		"00000000000000000000" &
		"101010000101000011" &
		"00000000000000000000" &
		"111000100101111010" &
		"00000000000000000000" &
		"111100010001011001" &
		"00000000000000000000" &
		"101101010011110" &
		"00000000000000000000" &
		"111111100100011111" &
		"00000000000000000000" &
		"00111110111001011" &
		"00000000000000000000" &
		"101100011010001111" &
		"00000000000000000000" &
		"011101011010100101" &
		"00000000000000000000" &
		"01100010001000010" &
		"00000000000000000000" &
		"001110111010010000" &
		"00000000000000000000" &
		"011111100101101111" &
		"00000000000000000000" &
		"0110101011000101" &
		"00000000000000000000" &
		"0010011010000110" &
		"00000000000000000000" &
		"011001001011010011" &
		"00000000000000000000" &
		"10110000010001101" &
		"00000000000000000000" &
		"001110110111010" &
		"00000000000000000000" &
		"001001100101111010" &
		"00000000000000000000" &
		"01101011100100110" &
		"00000000000000000000" &
		"01111100000000" &
		"00000000000000000000" &
		"101000011011111000" &
		"00000000000000000000" &
		"10110011101101101" &
		"00000000000000000000" &
		"1011100101011011" &
		"00000000000000000000" &
		"111110100101001001" &
		"00000000000000000000" &
		"001111001111100000" &
		"00000000000000000000" &
		"0010110100010010" &
		"00000000000000000000" &
		"011010111011000010" &
		"00000000000000000000" &
		"1010111111010101" &
		"00000000000000000000" &
		"0011101001101" &
		"00000000000000000000" &
		"111011000100110111" &
		"00000000000000000000" &
		"001000000111010001" &
		"00000000000000000000" &
		"10100110000011110" &
		"00000000000000000000" &
		"011101100000100010" &
		"00000000000000000000" &
		"00111011100001111" &
		"00000000000000000000" &
		"1111001000111101" &
		"00000000000000000000" &
		"10100011010011100" &
		"00000000000000000000" &
		"001001010100100011" &
		"00000000000000000000" &
		"001010111101011000" &
		"00000000000000000000" &
		"001100001101000000" &
		"00000000000000000000" &
		"01110000001101" &
		"00000000000000000000" &
		"111111011101101000" &
		"00000000000000000000" &
		"00101100001111000" &
		"00000000000000000000" &
		"1111111111101100" &
		"00000000000000000000" &
		"0111000101001000" &
		"00000000000000000000" &
		"001111110100111111" &
		"00000000000000000000" &
		"001110011101000111" &
		"00000000000000000000" &
		"001000111100010" &
		"00000000000000000000" &
		"0010011011010000" &
		"00000000000000000000" &
		"011000111110100" &
		"00000000000000000000" &
		"001101011111001010" &
		"00000000000000000000" &
		"01110111000110010" &
		"00000000000000000000" &
		"10100010101100000" &
		"00000000000000000000" &
		"101101110001010100" &
		"00000000000000000000" &
		"101011100001000110" &
		"00000000000000000000" &
		"00100001000100010" &
		"00000000000000000000" &
		"001111101000010000" &
		"00000000000000000000" &
		"011110000111100011" &
		"00000000000000000000" &
		"10111101101100111" &
		"00000000000000000000" &
		"11110000010100101" &
		"00000000000000000000" &
		"101011011001000110" &
		"00000000000000000000" &
		"001101000100011100" &
		"00000000000000000000" &
		"011001111000100" &
		"00000000000000000000" &
		"1111110001000011" &
		"00000000000000000000" &
		"011111000100011000" &
		"00000000000000000000" &
		"001000100110000010" &
		"00000000000000000000" &
		"101111100001100110" &
		"00000000000000000000" &
		"011011010011010000" &
		"00000000000000000000" &
		"111001101100100" &
		"00000000000000000000" &
		"011011111001000000" &
		"00000000000000000000" &
		"111110111100110001" &
		"00000000000000000000" &
		"101111000111101111" &
		"00000000000000000000" &
		"10100111100000010" &
		"00000000000000000000" &
		"01111010010111" &
		"00000000000000000000" &
		"10100001110010010" &
		"00000000000000000000" &
		"001100001110101100" &
		"00000000000000000000" &
		"00101101111000110" &
		"00000000000000000000" &
		"01111010000010" &
		"00000000000000000000" &
		"111011101101001011" &
		"00000000000000000000" &
		"101100111110001000" &
		"00000000000000000000" &
		"111000110010010101" &
		"00000000000000000000" &
		"01100000001101111" &
		"00000000000000000000" &
		"10101010110010000" &
		"00000000000000000000" &
		"10111000001111111" &
		"00000000000000000000" &
		"001100111010" &
		"00000000000000000000" &
		"1110110110110011" &
		"00000000000000000000" &
		"011100000000111000" &
		"00000000000000000000" &
		"111101101000110110" &
		"00000000000000000000" &
		"0110010001010100" &
		"00000000000000000000" &
		"001110111101100" &
		"00000000000000000000" &
		"011001110101010001" &
		"00000000000000000000" &
		"11111001101010011" &
		"00000000000000000000" &
		"001001011000111110" &
		"00000000000000000000" &
		"101110100000010101" &
		"00000000000000000000" &
		"01111100010110001" &
		"00000000000000000000" &
		"101000010100100001" &
		"00000000000000000000" &
		"00111101110001101" &
		"00000000000000000000" &
		"1111000000100100" &
		"00000000000000000000" &
		"1010110111001010" &
		"00000000000000000000" &
		"1110100110110001" &
		"00000000000000000000" &
		"0010001001101000" &
		"00000000000000000000" &
		"001010010110101" &
		"00000000000000000000" &
		"0111101011111" &
		"00000000000000000000" &
		"1010101010100011" &
		"00000000000000000000" &
		"0110101001100001" &
		"00000000000000000000" &
		"0110001000001101" &
		"00000000000000000000" &
		"1010110001011110" &
		"00000000000000000000" &
		"101111000011100000" &
		"00000000000000000000" &
		"111110101001000101" &
		"00000000000000000000" &
		"001111100111000" &
		"00000000000000000000" &
		"011101011110000100" &
		"00000000000000000000" &
		"111001001111101" &
		"00000000000000000000" &
		"101101000100101101" &
		"00000000000000000000" &
		"0011001001111001" &
		"00000000000000000000" &
		"11101101001011001" &
		"00000000000000000000" &
		"001000100001011000" &
		"00000000000000000000" &
		"011011011000010011" &
		"00000000000000000000" &
		"111110001100111001" &
		"00000000000000000000" &
		"111111110001001110" &
		"00000000000000000000" &
		"00100010110110110" &
		"00000000000000000000" &
		"1010101100010100" &
		"00000000000000000000" &
		"10111010001010" &
		"00000000000000000000" &
		"11110010000101000" &
		"00000000000000000000" &
		"1110011000010100" &
		"00000000000000000000" &
		"001001000111100101" &
		"00000000000000000000" &
		"111000101101001011" &
		"00000000000000000000" &
		"011110110111000011" &
		"00000000000000000000" &
		"001010010100010001" &
		"00000000000000000000" &
		"00110000100100011" &
		"00000000000000000000" &
		"011010000111000110" &
		"00000000000000000000" &
		"001100110001101100" &
		"00000000000000000000" &
		"111101101010101110" &
		"00000000000000000000" &
		"01110000010010100" &
		"00000000000000000000" &
		"111110101100000101" &
		"00000000000000000000" &
		"111100101101001001" &
		"00000000000000000000" &
		"11110110011101011" &
		"00000000000000000000" &
		"11111010101111000" &
		"00000000000000000000" &
		"10100100111000110" &
		"00000000000000000000" &
		"111010001010011110" &
		"00000000000000000000" &
		"011000011001011010" &
		"00000000000000000000" &
		"00100111000001010" &
		"00000000000000000000" &
		"101010101001000101" &
		"00000000000000000000" &
		"00110101010110000" &
		"00000000000000000000" &
		"101011001110011111" &
		"00000000000000000000" &
		"0110010000101110" &
		"00000000000000000000" &
		"1111111100110001" &
		"00000000000000000000" &
		"10110101110110001" &
		"00000000000000000000" &
		"1010011010111010" &
		"00000000000000000000" &
		"1010111110001001" &
		"00000000000000000000" &
		"001010000011011111" &
		"00000000000000000000" &
		"1111000010100101" &
		"00000000000000000000" &
		"10101110001100100" &
		"00000000000000000000" &
		"11101100100011011" &
		"00000000000000000000" &
		"011001111100011010" &
		"00000000000000000000" &
		"101110111111111001" &
		"00000000000000000000" &
		"0110010110000111" &
		"00000000000000000000" &
		"101000011111010011" &
		"00000000000000000000" &
		"101101000010111011" &
		"00000000000000000000" &
		"01100000110100000" &
		"00000000000000000000" &
		"011101010001000011" &
		"00000000000000000000" &
		"00110101000010010" &
		"00000000000000000000" &
		"00111000011010010" &
		"00000000000000000000" &
		"10101001011010010" &
		"00000000000000000000" &
		"0010111110001" &
		"00000000000000000000" &
		"111111100010101" &
		"00000000000000000000" &
		"1011000101101001" &
		"00000000000000000000" &
		"111111001100001011" &
		"00000000000000000000" &
		"11101100000000000" &
		"00000000000000000000" &
		"11110110011110000" &
		"00000000000000000000" &
		"10110101000011110" &
		"00000000000000000000" &
		"011000101001001101" &
		"00000000000000000000" &
		"10100100101001100" &
		"00000000000000000000" &
		"111010011001100100" &
		"00000000000000000000" &
		"01101000101010010" &
		"00000000000000000000" &
		"111111101101001000" &
		"00000000000000000000" &
		"0011001100101001" &
		"00000000000000000000" &
		"111100100000011000" &
		"00000000000000000000" &
		"0111111101011000" &
		"00000000000000000000" &
		"101101111100101100" &
		"00000000000000000000" &
		"111110010001000" &
		"00000000000000000000" &
		"1011011000101010" &
		"00000000000000000000" &
		"011010000001010001" &
		"00000000000000000000" &
		"001111100001001110" &
		"00000000000000000000" &
		"0111011101011001" &
		"00000000000000000000" &
		"1011111010101100" &
		"00000000000000000000" &
		"11111011101111" &
		"00000000000000000000" &
		"001100010101011" &
		"00000000000000000000" &
		"101100101101" &
		"00000000000000000000" &
		"11110111101100111" &
		"00000000000000000000" &
		"101011101110111000" &
		"00000000000000000000" &
		"011111001000110011" &
		"00000000000000000000" &
		"00101101101011011" &
		"00000000000000000000" &
		"011001110001010011" &
		"00000000000000000000" &
		"0110100110110000" &
		"00000000000000000000" &
		"011110100110001001" &
		"00000000000000000000" &
		"001100100100000000" &
		"00000000000000000000" &
		"11111011101110001" &
		"00000000000000000000" &
		"11111001110100000" &
		"00000000000000000000" &
		"00101010111111111" &
		"00000000000000000000" &
		"011001101101000010" &
		"00000000000000000000" &
		"101100000110011010" &
		"00000000000000000000" &
		"00111111001110001" &
		"00000000000000000000" &
		"101011100110000010" &
		"00000000000000000000" &
		"111000101000101110" &
		"00000000000000000000" &
		"101110100110010100" &
		"00000000000000000000" &
		"001100110101111111" &
		"00000000000000000000" &
		"00111111011" &
		"00000000000000000000" &
		"011101111111001110" &
		"00000000000000000000" &
		"111000011000000101" &
		"00000000000000000000" &
		"101011111010111111" &
		"00000000000000000000" &
		"101110111110010100" &
		"00000000000000000000" &
		"001000100000101001" &
		"00000000000000000000" &
		"10101010101010100" &
		"00000000000000000000" &
		"011100000100111101" &
		"00000000000000000000" &
		"101101111000000111" &
		"00000000000000000000" &
		"11111001010110011" &
		"00000000000000000000" &
		"00100100101111001" &
		"00000000000000000000" &
		"00101000011011000" &
		"00000000000000000000" &
		"011010110001000010" &
		"00000000000000000000" &
		"01111011101100010" &
		"00000000000000000000" &
		"00111001101000101" &
		"00000000000000000000" &
		"011100111000010110" &
		"00000000000000000000" &
		"101001001110010110" &
		"00000000000000000000" &
		"111111000110011001" &
		"00000000000000000000" &
		"1110111000111111" &
		"00000000000000000000" &
		"011010010010111100" &
		"00000000000000000000" &
		"101000111100111001" &
		"00000000000000000000" &
		"101001011101010111" &
		"00000000000000000000" &
		"111100101110011111" &
		"00000000000000000000" &
		"01100010110001001" &
		"00000000000000000000" &
		"111011011000011111" &
		"00000000000000000000" &
		"11100011001100010" &
		"00000000000000000000" &
		"101011111110111001" &
		"00000000000000000000" &
		"111010101100010110" &
		"00000000000000000000" &
		"1010101101111000" &
		"00000000000000000000" &
		"1010001100111" &
		"00000000000000000000" &
		"1111001001000101" &
		"00000000000000000000" &
		"10110011110110" &
		"00000000000000000000" &
		"111100101111001101" &
		"00000000000000000000" &
		"001101100110001111" &
		"00000000000000000000" &
		"11100000000110010" &
		"00000000000000000000" &
		"111101100111101011" &
		"00000000000000000000" &
		"1110000001001" &
		"00000000000000000000" &
		"01101010001101001" &
		"00000000000000000000" &
		"10100110001101100" &
		"00000000000000000000" &
		"101101001010000010" &
		"00000000000000000000" &
		"001000101000011000" &
		"00000000000000000000" &
		"11100111000010101" &
		"00000000000000000000" &
		"001010000010001111" &
		"00000000000000000000" &
		"1011110100001110" &
		"00000000000000000000" &
		"0011100000111111" &
		"00000000000000000000" &
		"00110100110110000" &
		"00000000000000000000" &
		"101101110011101100" &
		"00000000000000000000" &
		"101010110100111111" &
		"00000000000000000000" &
		"001101011011110010" &
		"00000000000000000000" &
		"011100100111100" &
		"00000000000000000000" &
		"11110001010110111" &
		"00000000000000000000" &
		"111000100110011101" &
		"00000000000000000000" &
		"0110100111101000" &
		"00000000000000000000" &
		"011011001011101101" &
		"00000000000000000000" &
		"0110100000010111" &
		"00000000000000000000" &
		"111000011111001010" &
		"00000000000000000000" &
		"001101000100110100" &
		"00000000000000000000" &
		"101011001110111111" &
		"00000000000000000000" &
		"001110001111111010" &
		"00000000000000000000" &
		"0111000100110110" &
		"00000000000000000000" &
		"111100101111010000" &
		"00000000000000000000" &
		"10110011110000011" &
		"00000000000000000000" &
		"011111001100011101" &
		"00000000000000000000" &
		"10100110001010010" &
		"00000000000000000000" &
		"01111011100001001" &
		"00000000000000000000" &
		"10100110100010" &
		"00000000000000000000" &
		"001100100011100111" &
		"00000000000000000000" &
		"0111100111000010" &
		"00000000000000000000" &
		"1111100101101110" &
		"00000000000000000000" &
		"01100100100111110" &
		"00000000000000000000" &
		"01110111101111111" &
		"00000000000000000000" &
		"11111001111110101" &
		"00000000000000000000" &
		"111100100111100101" &
		"00000000000000000000" &
		"101001000011000101" &
		"00000000000000000000" &
		"101011100010010010" &
		"00000000000000000000" &
		"101100111101011011" &
		"00000000000000000000" &
		"001110110001100011" &
		"00000000000000000000" &
		"111101001010000111" &
		"00000000000000000000" &
		"111100000000101110" &
		"00000000000000000000" &
		"00111110100011001" &
		"00000000000000000000" &
		"011111011110011001" &
		"00000000000000000000" &
		"011010011000101110" &
		"00000000000000000000" &
		"00101011111" &
		"00000000000000000000" &
		"1010010110" &
		"00000000000000000000" &
		"00110010110100111" &
		"00000000000000000000" &
		"101010000110001000" &
		"00000000000000000000" &
		"1011011000010000" &
		"00000000000000000000" &
		"10110001000111" &
		"00000000000000000000" &
		"01110001110100100" &
		"00000000000000000000" &
		"0111000001010101" &
		"00000000000000000000" &
		"111110011000001010" &
		"00000000000000000000" &
		"10100111010110001" &
		"00000000000000000000" &
		"101000000111011111" &
		"00000000000000000000" &
		"111000001101111100" &
		"00000000000000000000" &
		"11110100110001010" &
		"00000000000000000000" &
		"10110111110000000" &
		"00000000000000000000" &
		"111001000001000" &
		"00000000000000000000" &
		"01110111010110100" &
		"00000000000000000000" &
		"101011101111010110" &
		"00000000000000000000" &
		"1111001001011010" &
		"00000000000000000000" &
		"101111110011010110" &
		"00000000000000000000" ;

    -- Channel 2 -> MEM[1] -> 162
    -- Channel 1 -> MEM[2] -> 75

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (
				11343 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				62792 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				758 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				22696 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				49296 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				10690 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				50259 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				40839 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				28805 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				47057 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				57736 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				31915 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				36892 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				33537 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				2798 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				30969 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				30480 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				15196 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				16503 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				42727 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				24620 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				3540 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				6843 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				14214 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				32430 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				1227 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				42584 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				22281 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				39371 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				59372 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				38443 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				16463 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				18099 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				4886 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				12803 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				53732 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				13559 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				25760 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				20871 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				16762 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				5520 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				2910 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				36362 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				50346 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				1295 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				36713 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				25771 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				89 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				21756 => STD_LOGIC_VECTOR(to_unsigned(131, 8)),
				32606 => STD_LOGIC_VECTOR(to_unsigned(4, 8)),
				52113 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				59278 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				30991 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				13348 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				37879 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				2457 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				29889 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				50307 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				56221 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				5490 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				26870 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				50427 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				37817 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				48753 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				15577 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				9772 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				23562 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				27049 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				25312 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				7631 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				15848 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				39825 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				2874 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				27164 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				13648 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				34003 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				26299 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				11419 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				59503 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				49068 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				59982 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				50553 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				28190 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				29912 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				48835 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				20837 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				7158 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				56520 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				62904 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				14040 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				35800 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				51511 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				50505 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				10146 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				33929 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				22120 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				63081 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				18540 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				29320 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				16855 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				19063 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				59462 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				7287 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				30374 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				35319 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				25337 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				59731 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				17351 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				55567 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				21101 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				47691 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				28895 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				33813 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				3087 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				38803 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				64947 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				18181 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				22782 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				1476 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				11391 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				1755 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				50816 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				55516 => STD_LOGIC_VECTOR(to_unsigned(36, 8)),
				2693 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				32165 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				21480 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				13256 => STD_LOGIC_VECTOR(to_unsigned(192, 8)),
				33448 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				63392 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				61358 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				64661 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				49825 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				14441 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				14419 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				34739 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				50454 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				13522 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				38574 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				793 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				20988 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				23534 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				42387 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				50412 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				54679 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				58223 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				44005 => STD_LOGIC_VECTOR(to_unsigned(198, 8)),
				47221 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				38456 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				63797 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				35342 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				19481 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				16154 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				33453 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				44222 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				51167 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				19271 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				33380 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				12606 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				24727 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				30578 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				53499 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				58183 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				44941 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				29552 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				35734 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				47975 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				16652 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				43342 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				50208 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				56514 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				9036 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				54431 => STD_LOGIC_VECTOR(to_unsigned(134, 8)),
				25589 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				36485 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				55913 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				59106 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				38073 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				41444 => STD_LOGIC_VECTOR(to_unsigned(173, 8)),
				52321 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				5236 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				15679 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				58330 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				15837 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				21501 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				28587 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				13647 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				18766 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				5091 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				62970 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				50538 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				50035 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				42263 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				17077 => STD_LOGIC_VECTOR(to_unsigned(93, 8)),
				29524 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				24470 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				43981 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				28817 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				46738 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				53235 => STD_LOGIC_VECTOR(to_unsigned(186, 8)),
				22670 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				11828 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				46253 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				56695 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				13948 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				1792 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				50123 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				26017 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				211 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				36309 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				27695 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				57570 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				60707 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				8337 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				15246 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				27757 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				30669 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				51854 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				36048 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				62073 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				49570 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				37660 => STD_LOGIC_VECTOR(to_unsigned(53, 8)),
				63978 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				55068 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				40674 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				37131 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				47978 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				17014 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				38632 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				43572 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				210 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				7011 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				57201 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				30904 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				816 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				20402 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				28608 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				28105 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				30412 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				52300 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				19653 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				44250 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				54789 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				62241 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				56044 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				64137 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				14703 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				63025 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				26750 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				20155 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				743 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				2770 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				40944 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				26707 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				13393 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				17058 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				11982 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				15060 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				57100 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				59474 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				42771 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				34397 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				51422 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				36092 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				15270 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				38549 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				63015 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				60422 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				19929 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				17387 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				44558 => STD_LOGIC_VECTOR(to_unsigned(19, 8)),
				18884 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				54696 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				56084 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				40439 => STD_LOGIC_VECTOR(to_unsigned(150, 8)),
				52662 => STD_LOGIC_VECTOR(to_unsigned(145, 8)),
				4729 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				11151 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				13005 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				31384 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				50880 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				19974 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				16096 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				48435 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				7367 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				20376 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				2951 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				45737 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				24190 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				38824 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				42403 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				47312 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				40545 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				33293 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				43175 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				28108 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				731 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				41752 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				18414 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				6837 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				16079 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				57554 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				62396 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				3529 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				12664 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				36772 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				60255 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				2727 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				26687 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				47529 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				55200 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				30821 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				52664 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				49471 => STD_LOGIC_VECTOR(to_unsigned(194, 8)),
				51914 => STD_LOGIC_VECTOR(to_unsigned(73, 8)),
				54148 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				8498 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				47910 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				7294 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				35077 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				9362 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				32864 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				36858 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				57860 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				33809 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				55677 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				49267 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				58936 => STD_LOGIC_VECTOR(to_unsigned(29, 8)),
				6078 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				51249 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				48819 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				54537 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				51796 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				17967 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				51203 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				22529 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				21848 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				10895 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				38505 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				4611 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				31104 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				8794 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				24350 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				14108 => STD_LOGIC_VECTOR(to_unsigned(237, 8)),
				22959 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				17777 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				57614 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				54842 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				47696 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				55205 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				37701 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				24504 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				43217 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				26792 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				61765 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				56965 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				57636 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				16839 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				46190 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				33155 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				52335 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				42954 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				13555 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				35221 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				6358 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				64466 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				31340 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				58650 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				10954 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				59398 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				22683 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				56532 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				11355 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				24563 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				39605 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				20091 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				30321 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				44610 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				28816 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				60644 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				6269 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				48446 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				54241 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				9185 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				61587 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				46944 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				23696 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				47038 => STD_LOGIC_VECTOR(to_unsigned(80, 8)),
				39817 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				882 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				9768 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				18408 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				58939 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				26598 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				5365 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				39298 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				16465 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				57097 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				1084 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				44574 => STD_LOGIC_VECTOR(to_unsigned(117, 8)),
				46 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				46738 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				17970 => STD_LOGIC_VECTOR(to_unsigned(136, 8)),
				38681 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				63720 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				43649 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				14598 => STD_LOGIC_VECTOR(to_unsigned(209, 8)),
				27146 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				31499 => STD_LOGIC_VECTOR(to_unsigned(84, 8)),
				11688 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				6800 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				64511 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				61718 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				43166 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				34021 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				54106 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				58940 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				25686 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				25020 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				39369 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				61946 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				27748 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				40716 => STD_LOGIC_VECTOR(to_unsigned(231, 8)),
				3120 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				58360 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				52428 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				35078 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				29401 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				28349 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				64686 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				31224 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				6408 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				14661 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				17163 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				4813 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				7929 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				60587 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				22002 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				59950 => STD_LOGIC_VECTOR(to_unsigned(42, 8)),
				25512 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				58511 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				20670 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				17541 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				38764 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				33627 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				61121 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				31424 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				56141 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				44108 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				31469 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				9226 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				2635 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				31715 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				35925 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				8092 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				53526 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				36085 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				27502 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				507 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				46752 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				18809 => STD_LOGIC_VECTOR(to_unsigned(184, 8)),
				20848 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				18940 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				28039 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				10775 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				43979 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				40295 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				3864 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				39389 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				48143 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				35608 => STD_LOGIC_VECTOR(to_unsigned(210, 8)),
				49675 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				60222 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				749 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				5351 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				3468 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				9853 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				64335 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				26072 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				51176 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				50954 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				53076 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				2726 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				55225 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				13106 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				19776 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				33916 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				59438 => STD_LOGIC_VECTOR(to_unsigned(90, 8)),
				61555 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				4132 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				4341 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				21590 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				25377 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				63440 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				52646 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				27759 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				60476 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				44203 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				56478 => STD_LOGIC_VECTOR(to_unsigned(188, 8)),
				35221 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				4714 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				55347 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				8381 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				44840 => STD_LOGIC_VECTOR(to_unsigned(215, 8)),
				48693 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				44888 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				60131 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				43141 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				45968 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				52834 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				58992 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				59646 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				26989 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				31521 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				36953 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				13493 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				14070 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				54262 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				43665 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				11374 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				29115 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				60681 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				47406 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				8305 => STD_LOGIC_VECTOR(to_unsigned(155, 8)),
				31928 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				24312 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				24808 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				10096 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				46352 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				58627 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				30783 => STD_LOGIC_VECTOR(to_unsigned(30, 8)),
				42305 => STD_LOGIC_VECTOR(to_unsigned(180, 8)),
				20634 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				3781 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				55542 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				64778 => STD_LOGIC_VECTOR(to_unsigned(235, 8)),
				51188 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				39723 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				48304 => STD_LOGIC_VECTOR(to_unsigned(32, 8)),
				46083 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				31980 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				60902 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				5401 => STD_LOGIC_VECTOR(to_unsigned(225, 8)),
				12549 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				63610 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				12902 => STD_LOGIC_VECTOR(to_unsigned(0, 8)),
				63887 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				41960 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				31725 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				14946 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				59629 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				40853 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				40894 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				13803 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				44060 => STD_LOGIC_VECTOR(to_unsigned(170, 8)),
				44059 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				12714 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				12585 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				36309 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				64535 => STD_LOGIC_VECTOR(to_unsigned(217, 8)),
				33199 => STD_LOGIC_VECTOR(to_unsigned(174, 8)),
				3972 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				40847 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				31454 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				10483 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				21772 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				63488 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				3852 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				64251 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				10782 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				30552 => STD_LOGIC_VECTOR(to_unsigned(139, 8)),
				43625 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				26581 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				38599 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				25806 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				40060 => STD_LOGIC_VECTOR(to_unsigned(189, 8)),
				8678 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				13221 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				31385 => STD_LOGIC_VECTOR(to_unsigned(253, 8)),
				5904 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				10293 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				58449 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				22431 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				20849 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				57700 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				59199 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				46633 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				42483 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				52214 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				11811 => STD_LOGIC_VECTOR(to_unsigned(246, 8)),
				12247 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				709 => STD_LOGIC_VECTOR(to_unsigned(51, 8)),
				61847 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				50483 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				28821 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				64429 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				27053 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				51371 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				37882 => STD_LOGIC_VECTOR(to_unsigned(214, 8)),
				5058 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				34574 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				20693 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				6095 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				52716 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				38887 => STD_LOGIC_VECTOR(to_unsigned(130, 8)),
				61930 => STD_LOGIC_VECTOR(to_unsigned(140, 8)),
				44255 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				51857 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				28746 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				2511 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				15325 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				55859 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				22220 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				53852 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				55788 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				43603 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				34050 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				7704 => STD_LOGIC_VECTOR(to_unsigned(166, 8)),
				27297 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				652 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				39324 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				60815 => STD_LOGIC_VECTOR(to_unsigned(48, 8)),
				43386 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				55120 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				57257 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				55595 => STD_LOGIC_VECTOR(to_unsigned(203, 8)),
				63143 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				22452 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				47617 => STD_LOGIC_VECTOR(to_unsigned(156, 8)),
				61706 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				10943 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				9424 => STD_LOGIC_VECTOR(to_unsigned(33, 8)),
				4398 => STD_LOGIC_VECTOR(to_unsigned(222, 8)),
				27218 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				41957 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				7477 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				58266 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				18043 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				36106 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				25848 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				48453 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				35734 => STD_LOGIC_VECTOR(to_unsigned(1, 8)),
				7504 => STD_LOGIC_VECTOR(to_unsigned(193, 8)),
				50296 => STD_LOGIC_VECTOR(to_unsigned(12, 8)),
				46132 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				62524 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				44098 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				38211 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				46201 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				61864 => STD_LOGIC_VECTOR(to_unsigned(106, 8)),
				36336 => STD_LOGIC_VECTOR(to_unsigned(8, 8)),
				8526 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				26720 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				48293 => STD_LOGIC_VECTOR(to_unsigned(245, 8)),
				14235 => STD_LOGIC_VECTOR(to_unsigned(152, 8)),
				1577 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				34545 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				18744 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				46243 => STD_LOGIC_VECTOR(to_unsigned(146, 8)),
				59407 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				14269 => STD_LOGIC_VECTOR(to_unsigned(46, 8)),
				21711 => STD_LOGIC_VECTOR(to_unsigned(35, 8)),
				28282 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				17180 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				11296 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				64046 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				27440 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				10553 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				26615 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				49586 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				26602 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				63903 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				30154 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				50271 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				47284 => STD_LOGIC_VECTOR(to_unsigned(172, 8)),
				6069 => STD_LOGIC_VECTOR(to_unsigned(249, 8)),
				28531 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				40093 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				20065 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				39559 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				6641 => STD_LOGIC_VECTOR(to_unsigned(62, 8)),
				18459 => STD_LOGIC_VECTOR(to_unsigned(49, 8)),
				8855 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				28347 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				20387 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				5609 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				53249 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				21808 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				32597 => STD_LOGIC_VECTOR(to_unsigned(242, 8)),
				47159 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				29949 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				44795 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				21921 => STD_LOGIC_VECTOR(to_unsigned(65, 8)),
				62339 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				32865 => STD_LOGIC_VECTOR(to_unsigned(114, 8)),
				46724 => STD_LOGIC_VECTOR(to_unsigned(236, 8)),
				41283 => STD_LOGIC_VECTOR(to_unsigned(229, 8)),
				35194 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				50265 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				6814 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				63775 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				32203 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				50831 => STD_LOGIC_VECTOR(to_unsigned(197, 8)),
				54949 => STD_LOGIC_VECTOR(to_unsigned(99, 8)),
				17474 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				61072 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				63855 => STD_LOGIC_VECTOR(to_unsigned(3, 8)),
				10949 => STD_LOGIC_VECTOR(to_unsigned(141, 8)),
				9862 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				37587 => STD_LOGIC_VECTOR(to_unsigned(118, 8)),
				24717 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				7610 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				39290 => STD_LOGIC_VECTOR(to_unsigned(232, 8)),
				22310 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				3840 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				34552 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				26477 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				14683 => STD_LOGIC_VECTOR(to_unsigned(228, 8)),
				59721 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				62432 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				11538 => STD_LOGIC_VECTOR(to_unsigned(120, 8)),
				44738 => STD_LOGIC_VECTOR(to_unsigned(221, 8)),
				12245 => STD_LOGIC_VECTOR(to_unsigned(165, 8)),
				1869 => STD_LOGIC_VECTOR(to_unsigned(56, 8)),
				45367 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				33233 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				19486 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				55330 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				30479 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				12861 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				18076 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				38179 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				44888 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				49984 => STD_LOGIC_VECTOR(to_unsigned(47, 8)),
				3085 => STD_LOGIC_VECTOR(to_unsigned(39, 8)),
				63336 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				22648 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				16364 => STD_LOGIC_VECTOR(to_unsigned(126, 8)),
				12616 => STD_LOGIC_VECTOR(to_unsigned(219, 8)),
				64831 => STD_LOGIC_VECTOR(to_unsigned(10, 8)),
				59207 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				4578 => STD_LOGIC_VECTOR(to_unsigned(67, 8)),
				9936 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				4596 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				55242 => STD_LOGIC_VECTOR(to_unsigned(227, 8)),
				28210 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				17760 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				56404 => STD_LOGIC_VECTOR(to_unsigned(199, 8)),
				47174 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				16930 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				64016 => STD_LOGIC_VECTOR(to_unsigned(181, 8)),
				57827 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				31591 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				24741 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				46662 => STD_LOGIC_VECTOR(to_unsigned(204, 8)),
				53532 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				5060 => STD_LOGIC_VECTOR(to_unsigned(142, 8)),
				15427 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				61720 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				35202 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				63590 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				46288 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				4964 => STD_LOGIC_VECTOR(to_unsigned(175, 8)),
				48704 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				61233 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				61935 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				20226 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				3735 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				17298 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				50092 => STD_LOGIC_VECTOR(to_unsigned(100, 8)),
				23494 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				3714 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				47947 => STD_LOGIC_VECTOR(to_unsigned(27, 8)),
				53128 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				35989 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				16495 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				21904 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				28799 => STD_LOGIC_VECTOR(to_unsigned(119, 8)),
				826 => STD_LOGIC_VECTOR(to_unsigned(89, 8)),
				11699 => STD_LOGIC_VECTOR(to_unsigned(147, 8)),
				49208 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				55862 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				9300 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				7660 => STD_LOGIC_VECTOR(to_unsigned(163, 8)),
				40273 => STD_LOGIC_VECTOR(to_unsigned(247, 8)),
				29523 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				38462 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				59413 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				30897 => STD_LOGIC_VECTOR(to_unsigned(21, 8)),
				34081 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				31629 => STD_LOGIC_VECTOR(to_unsigned(148, 8)),
				12324 => STD_LOGIC_VECTOR(to_unsigned(205, 8)),
				11722 => STD_LOGIC_VECTOR(to_unsigned(64, 8)),
				10673 => STD_LOGIC_VECTOR(to_unsigned(76, 8)),
				8808 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				5301 => STD_LOGIC_VECTOR(to_unsigned(220, 8)),
				1887 => STD_LOGIC_VECTOR(to_unsigned(66, 8)),
				10915 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				10849 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				8717 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				11358 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				61664 => STD_LOGIC_VECTOR(to_unsigned(233, 8)),
				59973 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				7992 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				55172 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				4733 => STD_LOGIC_VECTOR(to_unsigned(161, 8)),
				53549 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				12921 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				23129 => STD_LOGIC_VECTOR(to_unsigned(252, 8)),
				34904 => STD_LOGIC_VECTOR(to_unsigned(52, 8)),
				46611 => STD_LOGIC_VECTOR(to_unsigned(96, 8)),
				58169 => STD_LOGIC_VECTOR(to_unsigned(71, 8)),
				64590 => STD_LOGIC_VECTOR(to_unsigned(208, 8)),
				17846 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				11028 => STD_LOGIC_VECTOR(to_unsigned(182, 8)),
				3722 => STD_LOGIC_VECTOR(to_unsigned(79, 8)),
				25640 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				9748 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				37349 => STD_LOGIC_VECTOR(to_unsigned(74, 8)),
				35659 => STD_LOGIC_VECTOR(to_unsigned(108, 8)),
				60867 => STD_LOGIC_VECTOR(to_unsigned(211, 8)),
				42257 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				24867 => STD_LOGIC_VECTOR(to_unsigned(6, 8)),
				41414 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				52332 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				55982 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				24724 => STD_LOGIC_VECTOR(to_unsigned(129, 8)),
				60165 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				52041 => STD_LOGIC_VECTOR(to_unsigned(31, 8)),
				27883 => STD_LOGIC_VECTOR(to_unsigned(116, 8)),
				30072 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				18886 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				41630 => STD_LOGIC_VECTOR(to_unsigned(102, 8)),
				34394 => STD_LOGIC_VECTOR(to_unsigned(57, 8)),
				19978 => STD_LOGIC_VECTOR(to_unsigned(91, 8)),
				43589 => STD_LOGIC_VECTOR(to_unsigned(135, 8)),
				27312 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				45983 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				9262 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				16177 => STD_LOGIC_VECTOR(to_unsigned(75, 8)),
				27569 => STD_LOGIC_VECTOR(to_unsigned(240, 8)),
				9914 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				12169 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				41183 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				12453 => STD_LOGIC_VECTOR(to_unsigned(38, 8)),
				23652 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				22811 => STD_LOGIC_VECTOR(to_unsigned(187, 8)),
				40730 => STD_LOGIC_VECTOR(to_unsigned(143, 8)),
				61433 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				9607 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				34771 => STD_LOGIC_VECTOR(to_unsigned(95, 8)),
				53435 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				16800 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				54339 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				27154 => STD_LOGIC_VECTOR(to_unsigned(241, 8)),
				28882 => STD_LOGIC_VECTOR(to_unsigned(83, 8)),
				21202 => STD_LOGIC_VECTOR(to_unsigned(254, 8)),
				1521 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				7957 => STD_LOGIC_VECTOR(to_unsigned(92, 8)),
				12649 => STD_LOGIC_VECTOR(to_unsigned(125, 8)),
				62219 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				22528 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				27888 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				27166 => STD_LOGIC_VECTOR(to_unsigned(34, 8)),
				35405 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				18764 => STD_LOGIC_VECTOR(to_unsigned(17, 8)),
				42596 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				20818 => STD_LOGIC_VECTOR(to_unsigned(201, 8)),
				64328 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				13097 => STD_LOGIC_VECTOR(to_unsigned(195, 8)),
				51224 => STD_LOGIC_VECTOR(to_unsigned(13, 8)),
				16216 => STD_LOGIC_VECTOR(to_unsigned(202, 8)),
				57132 => STD_LOGIC_VECTOR(to_unsigned(224, 8)),
				7304 => STD_LOGIC_VECTOR(to_unsigned(133, 8)),
				13866 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				41041 => STD_LOGIC_VECTOR(to_unsigned(138, 8)),
				63566 => STD_LOGIC_VECTOR(to_unsigned(97, 8)),
				14169 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				16044 => STD_LOGIC_VECTOR(to_unsigned(149, 8)),
				3823 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				6315 => STD_LOGIC_VECTOR(to_unsigned(37, 8)),
				813 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				28519 => STD_LOGIC_VECTOR(to_unsigned(86, 8)),
				48056 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				62003 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				23387 => STD_LOGIC_VECTOR(to_unsigned(177, 8)),
				40019 => STD_LOGIC_VECTOR(to_unsigned(55, 8)),
				10672 => STD_LOGIC_VECTOR(to_unsigned(238, 8)),
				59785 => STD_LOGIC_VECTOR(to_unsigned(196, 8)),
				51456 => STD_LOGIC_VECTOR(to_unsigned(70, 8)),
				30577 => STD_LOGIC_VECTOR(to_unsigned(212, 8)),
				29600 => STD_LOGIC_VECTOR(to_unsigned(144, 8)),
				22015 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				39746 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				49562 => STD_LOGIC_VECTOR(to_unsigned(101, 8)),
				32369 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				47490 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				35374 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				59796 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),
				52607 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				507 => STD_LOGIC_VECTOR(to_unsigned(88, 8)),
				57294 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				34309 => STD_LOGIC_VECTOR(to_unsigned(132, 8)),
				48831 => STD_LOGIC_VECTOR(to_unsigned(41, 8)),
				61332 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				34857 => STD_LOGIC_VECTOR(to_unsigned(239, 8)),
				21844 => STD_LOGIC_VECTOR(to_unsigned(20, 8)),
				49469 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				56839 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				29363 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
				18809 => STD_LOGIC_VECTOR(to_unsigned(16, 8)),
				20696 => STD_LOGIC_VECTOR(to_unsigned(14, 8)),
				44098 => STD_LOGIC_VECTOR(to_unsigned(68, 8)),
				30562 => STD_LOGIC_VECTOR(to_unsigned(124, 8)),
				29509 => STD_LOGIC_VECTOR(to_unsigned(158, 8)),
				52758 => STD_LOGIC_VECTOR(to_unsigned(103, 8)),
				37782 => STD_LOGIC_VECTOR(to_unsigned(40, 8)),
				61849 => STD_LOGIC_VECTOR(to_unsigned(112, 8)),
				11839 => STD_LOGIC_VECTOR(to_unsigned(59, 8)),
				42172 => STD_LOGIC_VECTOR(to_unsigned(123, 8)),
				36665 => STD_LOGIC_VECTOR(to_unsigned(234, 8)),
				38743 => STD_LOGIC_VECTOR(to_unsigned(105, 8)),
				52127 => STD_LOGIC_VECTOR(to_unsigned(216, 8)),
				17801 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				46623 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				18018 => STD_LOGIC_VECTOR(to_unsigned(15, 8)),
				49081 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				43798 => STD_LOGIC_VECTOR(to_unsigned(153, 8)),
				11128 => STD_LOGIC_VECTOR(to_unsigned(94, 8)),
				1127 => STD_LOGIC_VECTOR(to_unsigned(111, 8)),
				12869 => STD_LOGIC_VECTOR(to_unsigned(250, 8)),
				3318 => STD_LOGIC_VECTOR(to_unsigned(61, 8)),
				52173 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				55695 => STD_LOGIC_VECTOR(to_unsigned(121, 8)),
				16434 => STD_LOGIC_VECTOR(to_unsigned(191, 8)),
				55787 => STD_LOGIC_VECTOR(to_unsigned(60, 8)),
				1033 => STD_LOGIC_VECTOR(to_unsigned(54, 8)),
				21609 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				19564 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				53890 => STD_LOGIC_VECTOR(to_unsigned(169, 8)),
				35352 => STD_LOGIC_VECTOR(to_unsigned(157, 8)),
				19989 => STD_LOGIC_VECTOR(to_unsigned(244, 8)),
				41103 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				15630 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				14399 => STD_LOGIC_VECTOR(to_unsigned(168, 8)),
				27056 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				56556 => STD_LOGIC_VECTOR(to_unsigned(137, 8)),
				44351 => STD_LOGIC_VECTOR(to_unsigned(104, 8)),
				55026 => STD_LOGIC_VECTOR(to_unsigned(183, 8)),
				6460 => STD_LOGIC_VECTOR(to_unsigned(176, 8)),
				25271 => STD_LOGIC_VECTOR(to_unsigned(2, 8)),
				35229 => STD_LOGIC_VECTOR(to_unsigned(58, 8)),
				10728 => STD_LOGIC_VECTOR(to_unsigned(85, 8)),
				45805 => STD_LOGIC_VECTOR(to_unsigned(213, 8)),
				10263 => STD_LOGIC_VECTOR(to_unsigned(107, 8)),
				34762 => STD_LOGIC_VECTOR(to_unsigned(7, 8)),
				53556 => STD_LOGIC_VECTOR(to_unsigned(72, 8)),
				46015 => STD_LOGIC_VECTOR(to_unsigned(207, 8)),
				58362 => STD_LOGIC_VECTOR(to_unsigned(87, 8)),
				12598 => STD_LOGIC_VECTOR(to_unsigned(248, 8)),
				52176 => STD_LOGIC_VECTOR(to_unsigned(98, 8)),
				26499 => STD_LOGIC_VECTOR(to_unsigned(164, 8)),
				62237 => STD_LOGIC_VECTOR(to_unsigned(167, 8)),
				19538 => STD_LOGIC_VECTOR(to_unsigned(226, 8)),
				30473 => STD_LOGIC_VECTOR(to_unsigned(159, 8)),
				2466 => STD_LOGIC_VECTOR(to_unsigned(171, 8)),
				51431 => STD_LOGIC_VECTOR(to_unsigned(69, 8)),
				14786 => STD_LOGIC_VECTOR(to_unsigned(113, 8)),
				14702 => STD_LOGIC_VECTOR(to_unsigned(24, 8)),
				18750 => STD_LOGIC_VECTOR(to_unsigned(122, 8)),
				28543 => STD_LOGIC_VECTOR(to_unsigned(78, 8)),
				29685 => STD_LOGIC_VECTOR(to_unsigned(179, 8)),
				51685 => STD_LOGIC_VECTOR(to_unsigned(45, 8)),
				37061 => STD_LOGIC_VECTOR(to_unsigned(110, 8)),
				47250 => STD_LOGIC_VECTOR(to_unsigned(22, 8)),
				53083 => STD_LOGIC_VECTOR(to_unsigned(251, 8)),
				60515 => STD_LOGIC_VECTOR(to_unsigned(81, 8)),
				53895 => STD_LOGIC_VECTOR(to_unsigned(243, 8)),
				49198 => STD_LOGIC_VECTOR(to_unsigned(11, 8)),
				32025 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				63385 => STD_LOGIC_VECTOR(to_unsigned(154, 8)),
				42542 => STD_LOGIC_VECTOR(to_unsigned(230, 8)),
				351 => STD_LOGIC_VECTOR(to_unsigned(23, 8)),
				150 => STD_LOGIC_VECTOR(to_unsigned(28, 8)),
				26023 => STD_LOGIC_VECTOR(to_unsigned(151, 8)),
				41352 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				13840 => STD_LOGIC_VECTOR(to_unsigned(128, 8)),
				3143 => STD_LOGIC_VECTOR(to_unsigned(63, 8)),
				25508 => STD_LOGIC_VECTOR(to_unsigned(44, 8)),
				12373 => STD_LOGIC_VECTOR(to_unsigned(178, 8)),
				58890 => STD_LOGIC_VECTOR(to_unsigned(185, 8)),
				20145 => STD_LOGIC_VECTOR(to_unsigned(127, 8)),
				33247 => STD_LOGIC_VECTOR(to_unsigned(115, 8)),
				33660 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				27018 => STD_LOGIC_VECTOR(to_unsigned(218, 8)),
				28544 => STD_LOGIC_VECTOR(to_unsigned(160, 8)),
				4616 => STD_LOGIC_VECTOR(to_unsigned(109, 8)),
				28340 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),
				48086 => STD_LOGIC_VECTOR(to_unsigned(25, 8)),
				12890 => STD_LOGIC_VECTOR(to_unsigned(206, 8)),
				64726 => STD_LOGIC_VECTOR(to_unsigned(82, 8)),

                              
                                
                                OTHERS => "00000000"-- (OTHERS => '0')
                            );
                    
    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
            END IF;
        END IF;
    END PROCESS;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";
        -- wait for 10000 ns;
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        WAIT UNTIL tb_start = '1';
        ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  0
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  0
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(242, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  242
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  0
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  0
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  123
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  118
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  228
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  175
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  129
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  175
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  175
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  175
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  188
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  41
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  41
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  225
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  225
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  225
        ASSERT tb_z1 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  246
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  225
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  73
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  132
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  250
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  250
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  250
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  250
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  221
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  128
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  34
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  89
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  226
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(131, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  131
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  201
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  18
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  170
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  18
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  154
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(4, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  4
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  26
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  26
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  51
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  51
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  152
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  217
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  184
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  113
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  184
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  113
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  250
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  250
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  233
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  161
        ASSERT tb_z3 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  233
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  233
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  82
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  82
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  155
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  155
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  95
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  127
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  127
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  35
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  35
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  35
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  114
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  237
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  205
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  109
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  109
        ASSERT tb_z1 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  240
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  109
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  117
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  52
        ASSERT tb_z2 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  192
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(134, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  134
        ASSERT tb_z2 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  192
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  192
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  192
        ASSERT tb_z3 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  194
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  194
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  194
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  194
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  215
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  215
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  215
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  215
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  37
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  115
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  63
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  192
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(192, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  192
        ASSERT tb_z1 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  241
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  167
        ASSERT tb_z1 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  241
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(36, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  36
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  167
        ASSERT tb_z1 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  241
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  241
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  6
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  29
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  126
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  126
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  72
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  81
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  186
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  188
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  188
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  66
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  69
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  198
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  198
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(198, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  198
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  125
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  216
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  8
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  8
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  8
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  219
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  226
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  0
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  42
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  132
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  63
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  63
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  25
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  26
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(134, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  134
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(134, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  134
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(134, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  134
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  87
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  181
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  182
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  102
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(173, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  173
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  125
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  194
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  125
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  125
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  177
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  155
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  79
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  249
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  79
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(186, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  186
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  191
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  191
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(93, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  93
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  65
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  18
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  120
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  96
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  97
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  18
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  103
        ASSERT tb_z1 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  116
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  103
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  189
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  138
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  231
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  156
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(53, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  53
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  81
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  139
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  81
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  33
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  81
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  184
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  81
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  86
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  81
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  86
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  157
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  1
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  19
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  19
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  226
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  214
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  13
        ASSERT tb_z3 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  210
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  210
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  227
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  210
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  227
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  3
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  40
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  103
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  133
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  195
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  86
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  107
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  95
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  95
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  218
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  218
        ASSERT tb_z2 = std_logic_vector(to_unsigned(19, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  19
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  218
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  218
        ASSERT tb_z2 = std_logic_vector(to_unsigned(150, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  150
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  218
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  154
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  39
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  235
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(145, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  145
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  176
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  124
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  163
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  118
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  204
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  132
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  65
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  17
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  60
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  73
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  8
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  111
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  197
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  111
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  111
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  126
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  126
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  222
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  58
        ASSERT tb_z1 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  194
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(73, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  73
        ASSERT tb_z1 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  194
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(194, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  194
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  247
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  248
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  44
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  214
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  44
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  214
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  214
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  214
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  183
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  214
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  217
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  217
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  217
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  245
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  101
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  82
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  239
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  82
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  51
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(29, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  29
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  241
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  112
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  225
        ASSERT tb_z3 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  46
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  225
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  91
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  91
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  249
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(237, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  237
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  160
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  202
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  32
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  238
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  205
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  127
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  127
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  133
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  181
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  149
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  76
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  159
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  64
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  159
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  108
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  143
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  108
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  94
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  94
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  94
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  222
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  94
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  58
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  139
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  182
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  182
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  182
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  239
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  172
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  214
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  238
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  221
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  221
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  75
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  208
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  80
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  124
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(80, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  80
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  127
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  127
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  117
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  183
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  117
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(117, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  117
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(136, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  136
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  203
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  187
        ASSERT tb_z2 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  144
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  187
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(209, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  209
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  189
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  180
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  157
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  221
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(84, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  84
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  253
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  103
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  225
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  39
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  120
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  10
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(231, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  231
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  230
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  24
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  24
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  174
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  174
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  174
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  142
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  67
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  118
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  67
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  118
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  101
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  75
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  8
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  8
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(42, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  42
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  8
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  8
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  82
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  133
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  82
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  147
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  82
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  147
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  147
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  35
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(146, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  146
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  35
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(146, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  146
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  70
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  70
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  0
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  66
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  66
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  23
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  139
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  250
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  180
        ASSERT tb_z1 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  250
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  250
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  163
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  163
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(184, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  184
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  163
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  228
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  228
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  203
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  112
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  62
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  112
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  62
        ASSERT tb_z1 = std_logic_vector(to_unsigned(210, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  210
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  157
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  62
        ASSERT tb_z1 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  232
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  157
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  62
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  157
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  199
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  157
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  199
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  199
        ASSERT tb_z1 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  109
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  199
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  166
        ASSERT tb_z1 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  121
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  166
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  166
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  25
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  25
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  25
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(90, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  90
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  21
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  15
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  166
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  106
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  208
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  208
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(188, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  188
        ASSERT tb_z1 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  232
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  232
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  128
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  140
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(215, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  215
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  15
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  205
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  205
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  196
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  227
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  141
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  105
        ASSERT tb_z1 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  108
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  105
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  40
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  13
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  167
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  48
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  156
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  135
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  156
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  92
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  193
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  207
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  12
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  12
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(155, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  155
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(30, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  30
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  75
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(235, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  235
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(180, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  180
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  97
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  152
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  35
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(32, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  32
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(225, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  225
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  24
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  24
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  0
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  14
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  246
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  18
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  211
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  211
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  101
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  211
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  20
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  211
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  144
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(170, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  170
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  217
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  217
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(217, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  217
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  56
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(174, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  174
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  148
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  148
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(139, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  139
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  208
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  159
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  193
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  105
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  113
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(253, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  253
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  25
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(189, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  189
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  54
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  38
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  38
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  38
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  167
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  74
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  201
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  22
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(246, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  246
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  158
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  81
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  205
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  205
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(51, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  51
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  229
        ASSERT tb_z2 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  221
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  221
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(214, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  214
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  245
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  140
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  138
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  14
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  130
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(130, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  130
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  46
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(140, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  140
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  46
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  92
        ASSERT tb_z1 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  46
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  46
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  82
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  211
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  82
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  126
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  126
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  7
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  207
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  118
        ASSERT tb_z1 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  179
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  118
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  118
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  49
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(166, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  166
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  27
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(203, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  203
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(48, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  48
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  244
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(156, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  156
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  213
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(33, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  33
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  83
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  10
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  78
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  12
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(222, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  222
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  183
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  87
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(1, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  1
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  149
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(193, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  193
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(12, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  12
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  179
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  91
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  157
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  100
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  59
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  22
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  8
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(8, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  8
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(245, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  245
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  199
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(106, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  106
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(152, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  152
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  22
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(146, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  146
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  165
        ASSERT tb_z1 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  110
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  110
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(35, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  35
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  199
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  61
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  49
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  228
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  109
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(46, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  46
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  105
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  254
        ASSERT tb_z1 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  6
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  6
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  6
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  6
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  6
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(249, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  249
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  244
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(172, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  172
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  244
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  49
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(49, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  49
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  126
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  252
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(62, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  62
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(242, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  242
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  121
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  25
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(65, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  65
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(114, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  114
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(229, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  229
        ASSERT tb_z3 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  148
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  148
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(236, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  236
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(99, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  99
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  57
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  92
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  92
        ASSERT tb_z1 = std_logic_vector(to_unsigned(3, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  3
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  92
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  202
        ASSERT tb_z1 = std_logic_vector(to_unsigned(141, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  141
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  202
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(197, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  197
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  202
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(118, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  118
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  239
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  126
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  11
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(232, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  232
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  34
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  220
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(228, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  228
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(120, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  120
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  56
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  113
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(56, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  56
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(165, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  165
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(221, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  221
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  206
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  164
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  206
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  239
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  206
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  178
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  204
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  47
        ASSERT tb_z1 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  27
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  47
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  178
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(47, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  47
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  85
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  26
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  85
        ASSERT tb_z1 = std_logic_vector(to_unsigned(39, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  39
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  85
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(10, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  10
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  135
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(67, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  67
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(219, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  219
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  54
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  38
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(199, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  199
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(227, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  227
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  82
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  119
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  76
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  133
        ASSERT tb_z3 = std_logic_vector(to_unsigned(126, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  126
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  133
        ASSERT tb_z3 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  163
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(181, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  181
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  163
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  23
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  163
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  142
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  163
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(142, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  142
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  9
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(204, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  204
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  28
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(175, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  175
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  178
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  21
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  135
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  27
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  233
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(100, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  100
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  187
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(27, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  27
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  233
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  108
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  79
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(147, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  147
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(89, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  89
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  163
        ASSERT tb_z1 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  111
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  163
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  177
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(163, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  163
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  137
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(119, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  119
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  137
        ASSERT tb_z1 = std_logic_vector(to_unsigned(247, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  247
        ASSERT tb_z2 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  116
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  137
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  116
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  137
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  224
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  16
        ASSERT tb_z3 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  205
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(205, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  205
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(148, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  148
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  238
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(21, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  21
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(64, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  64
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(66, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  66
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  38
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  40
        ASSERT tb_z2 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  216
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  40
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  40
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(76, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  76
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(220, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  220
        ASSERT tb_z1 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  40
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  40
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  248
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(233, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  233
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  240
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(161, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  161
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  41
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  52
        ASSERT tb_z1 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  243
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  52
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(252, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  252
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  52
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(71, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  71
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(52, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  52
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  251
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  129
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  251
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(182, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  182
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  251
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(208, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  208
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  251
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  251
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  44
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  74
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  44
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  74
        ASSERT tb_z1 = std_logic_vector(to_unsigned(96, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  96
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(74, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  74
        ASSERT tb_z1 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  211
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  11
        ASSERT tb_z1 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  211
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(211, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  211
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(6, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  6
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(108, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  108
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  151
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  110
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(31, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  31
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(116, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  116
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(79, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  79
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  124
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(129, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  129
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  218
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(91, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  91
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(135, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  135
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(57, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  57
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(102, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  102
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(240, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  240
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  185
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  122
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  122
        ASSERT tb_z3 = std_logic_vector(to_unsigned(75, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  75
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  122
        ASSERT tb_z3 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  38
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(38, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  38
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(143, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  143
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  69
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(95, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  95
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  16
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  112
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(241, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  241
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  83
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  97
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(83, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  83
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  254
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  254
        ASSERT tb_z3 = std_logic_vector(to_unsigned(187, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  187
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(254, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  254
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  125
        ASSERT tb_z3 = std_logic_vector(to_unsigned(92, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  92
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  125
        ASSERT tb_z3 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  68
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  125
        ASSERT tb_z3 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  123
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(125, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  125
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  34
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(34, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  34
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  17
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  104
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  224
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  234
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(201, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  201
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  13
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(17, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  17
        ASSERT tb_z3 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  13
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(13, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  13
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(224, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  224
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(202, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  202
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(195, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  195
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  97
        ASSERT tb_z1 = std_logic_vector(to_unsigned(138, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  138
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  97
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  70
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  97
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(133, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  133
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(97, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  97
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  37
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(149, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  149
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  37
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  37
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  37
        ASSERT tb_z1 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  88
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(37, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  37
        ASSERT tb_z1 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  60
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  60
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(55, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  55
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(238, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  238
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(177, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  177
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(86, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  86
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(212, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  212
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(70, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  70
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  44
        ASSERT tb_z1 = std_logic_vector(to_unsigned(196, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  196
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  44
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  230
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  44
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  248
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(101, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  101
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  248
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(144, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  144
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  248
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  248
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  18
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  7
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  63
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(41, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  41
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(88, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  88
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  151
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  20
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(132, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  132
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(239, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  239
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(16, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  16
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  158
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(68, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  68
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(14, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  14
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(124, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  124
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  9
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(18, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  18
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(112, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  112
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(103, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  103
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(40, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  40
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(234, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  234
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  105
        ASSERT tb_z3 = std_logic_vector(to_unsigned(59, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  59
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(123, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  123
        ASSERT tb_z2 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  105
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  105
        ASSERT tb_z3 = std_logic_vector(to_unsigned(216, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  216
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  105
        ASSERT tb_z3 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  110
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(105, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  105
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(15, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  15
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  153
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(94, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  94
        ASSERT tb_z3 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  153
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(153, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  153
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(111, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  111
        ASSERT tb_z3 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  250
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(250, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  250
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(158, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  158
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  213
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(191, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  191
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(60, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  60
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  169
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(61, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  61
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  168
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(121, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  121
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(54, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  54
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(157, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  157
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(169, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  169
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  78
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(168, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  168
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  127
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  213
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  127
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(137, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  137
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  127
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  176
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(244, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  244
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  176
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(2, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  2
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(176, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  176
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  58
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(85, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  85
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  58
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(213, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  213
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  58
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(58, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  58
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(183, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  183
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(104, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  104
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(72, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  72
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(107, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  107
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(7, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  7
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(207, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  207
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(248, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  248
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(164, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  164
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(167, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  167
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(226, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  226
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(87, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  87
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(159, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  159
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(98, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  98
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(113, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  113
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  24
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(122, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  122
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  24
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(24, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  24
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(179, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  179
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(171, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  171
        ASSERT tb_z3 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  45
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(110, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  110
        ASSERT tb_z3 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  45
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(22, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  22
        ASSERT tb_z3 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  45
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(69, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  69
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  45
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(45, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  45
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(243, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  243
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(81, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  81
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  28
        ASSERT tb_z1 = std_logic_vector(to_unsigned(78, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  78
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  28
        ASSERT tb_z1 = std_logic_vector(to_unsigned(154, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  154
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  28
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  23
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(251, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  251
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(23, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  23
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  28
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(28, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  28
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  25
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(128, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  128
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(230, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  230
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(44, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  44
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(11, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  11
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(63, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  63
        ASSERT tb_z3 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  185
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(127, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  127
        ASSERT tb_z3 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  185
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(185, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  185
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  160
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(115, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  115
        ASSERT tb_z3 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  218
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(218, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  218
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(178, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  178
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(160, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  160
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  25
        ASSERT tb_z3 = std_logic_vector(to_unsigned(109, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  109
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(25, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  25
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        WAIT UNTIL tb_done = '1';
        WAIT FOR CLOCK_PERIOD/2;

        ASSERT tb_z0 = std_logic_vector(to_unsigned(151, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure; --. Expected  151
        ASSERT tb_z1 = std_logic_vector(to_unsigned(9, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure; --. Expected  9
        ASSERT tb_z2 = std_logic_vector(to_unsigned(82, 8))  REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure; --. Expected  82
        ASSERT tb_z3 = std_logic_vector(to_unsigned(206, 8))  REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure; --. Expected  206
 
        
        ASSERT false REPORT "Simulation Ended! TEST PASSATO ()" SEVERITY failure;
    END PROCESS testRoutine;

END projecttb;
